/*
MIT License

Copyright (c) 2024 Elsie Rezinold Y

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
SOFTWARE.
*/
//`include "sixtyfourbit_lca.v"

module onetwoeightbit_lca (
    a,
    b,
    c,
    s
);


input [127:0] a,b;
input c;

output [127:0] s;
wire g1,p1;
wire g2,p2;

wire c2;

sixtyfourbit_lca uut_0 (
    a[63:0],
    b[63:0],
    c,
    s[63:0],
    g1,
    p1
);


assign c2 = g1 |(p1&c);

sixtyfourbit_lca uut_1 (
    a[127:64],
    b[127:64],
    c2,
    s[127:64],
    g2,
    p2
);


endmodule