/*
MIT License

Copyright (c) 2024 Elsie Rezinold Y

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
SOFTWARE.
*/
`define TAG 63:16
`define INDEX 15:6
`define OFFSET 5:0
module mem_cache (
clk,
rst_n,
i_cpu_address,  
i_cpu_din,
i_rd_valid,
i_wr_valid,          
o_cpu_dout_valid,
o_cpu_dout_data,
o_cache_busy,
miss,
o_mem_wr_data,
o_mem_rd_address,
o_mem_rd_valid,
o_mem_wr_address,
o_mem_wr_valid,
i_mem_rd_data,
i_mem_rd_data_valid,
i_mem_rd_data_tag,
cache_rd_wr_done,
mem_rd_wr_done
//valid_1,
//cache_mem_1,
//tag_1
);

parameter AWIDTH = 64, WIDTH=64,TAG_WIDTH=47;
input               clk;
input               rst_n;


input [AWIDTH-1:0]  i_cpu_address;  
input [WIDTH-1:0]              i_cpu_din;
input               i_rd_valid;
input               i_wr_valid;  
output reg          o_cpu_dout_valid;
output reg [WIDTH-1:0]  o_cpu_dout_data;
output reg              o_cache_busy;
output reg [WIDTH-1:0]  o_mem_wr_data;
output [AWIDTH-1:0] o_mem_rd_address;
output              o_mem_rd_valid;
output reg [AWIDTH-1:0] o_mem_wr_address;
output reg             o_mem_wr_valid;
input  [WIDTH-1:0]  i_mem_rd_data;
input               i_mem_rd_data_valid;
input  [AWIDTH-1:0] i_mem_rd_data_tag;
output              miss;
output reg cache_rd_wr_done;
output reg mem_rd_wr_done;
parameter CACHE_ACCESS=1'b0,MEM_ACCESS=1'b1;
reg  cs,ns;
//wire miss;
reg                        valid_1 [0:1023];
reg                        valid_2 [0:1023];
reg                    dirty_bit_1 [0:1023];
reg                    dirty_bit_2 [0:1023];
reg [TAG_WIDTH-1 :0]         tag_1 [0:1023];
reg [TAG_WIDTH-1 :0]         tag_2 [0:1023];
reg                  lru_counter_1 [0:1023];
reg                  lru_counter_2 [0:1023];
reg [WIDTH-1 :0]         cache_mem_1 [0:1023];
reg [WIDTH-1 :0]         cache_mem_2 [0:1023];
//reg cache_rd_wr_done;

always @(*) begin
  ns = 0;
  case(cs)
  CACHE_ACCESS: begin
    //if (!cache_rd_wr_done)
    if(miss)
      ns = MEM_ACCESS;
    else
      ns = CACHE_ACCESS;
  end
  MEM_ACCESS: begin
    if (mem_rd_wr_done)
      ns = CACHE_ACCESS;
    else
      ns = MEM_ACCESS;
  end
  endcase
end

always@(posedge clk or negedge rst_n)
  if(~rst_n)
    cs <= CACHE_ACCESS;
  else
    cs <= ns;

assign miss = ((i_rd_valid||i_wr_valid) &&!((valid_1[i_cpu_address[`INDEX]]&&(tag_1[i_cpu_address[`INDEX]]==i_cpu_address[`TAG]))|| (valid_2[i_cpu_address[`INDEX]]&&(tag_2[i_cpu_address[`INDEX]]==i_cpu_address[`TAG]))));

assign o_mem_rd_valid = miss;
assign o_mem_rd_address = i_cpu_address;

//assign o_cache_busy = !cache_rd_wr_done;

always@(posedge clk or negedge rst_n) begin
  if(rst_n) begin
    case(cs)
    CACHE_ACCESS : begin
      o_mem_wr_valid <= 0;
      mem_rd_wr_done <= 0;
      o_cache_busy   <= ((i_rd_valid||i_wr_valid) && !((valid_1[i_cpu_address[`INDEX]]&&(tag_1[i_cpu_address[`INDEX]]==i_cpu_address[`TAG])) || (valid_2[i_cpu_address[`INDEX]]&&(tag_2[i_cpu_address[`INDEX]]==i_cpu_address[`TAG]))));
      if(valid_1[i_cpu_address[`INDEX]]&&(tag_1[i_cpu_address[`INDEX]]==i_cpu_address[`TAG])) begin
        if(i_rd_valid) begin
          o_cpu_dout_valid <= i_rd_valid;
          o_cpu_dout_data  <= cache_mem_1[i_cpu_address[`INDEX]];
          lru_counter_1[i_cpu_address[`INDEX]] <= 1;
          lru_counter_2[i_cpu_address[`INDEX]] <= 0;
          cache_rd_wr_done                     <= 1;
        end
        else if(i_wr_valid) begin
          cache_mem_1[i_cpu_address[`INDEX]]   <= i_cpu_din;
          dirty_bit_1[i_cpu_address[`INDEX]]   <= 1'b1;
          tag_1[i_cpu_address[`INDEX]]         <= i_cpu_address[`TAG];
          lru_counter_1[i_cpu_address[`INDEX]] <= 1;
          lru_counter_2[i_cpu_address[`INDEX]] <= 0;
          cache_rd_wr_done <= 1;
        end                       
      end
      else if(valid_2[i_cpu_address[`INDEX]]&&(tag_2[i_cpu_address[`INDEX]]==i_cpu_address[`TAG])) begin
        if(i_wr_valid) begin
          cache_mem_2[i_cpu_address[`INDEX]]   <= i_cpu_din;
          dirty_bit_2[i_cpu_address[`INDEX]]   <= 1'b1;
          tag_2[i_cpu_address[`INDEX]]         <= i_cpu_address[`TAG];
          lru_counter_1[i_cpu_address[`INDEX]] <= 0;
          lru_counter_2[i_cpu_address[`INDEX]] <= 1;
          cache_rd_wr_done <= 1;
        end
        else if(i_rd_valid) begin
          o_cpu_dout_valid <= i_rd_valid;
          o_cpu_dout_data  <= cache_mem_2[i_cpu_address[`INDEX]];
          lru_counter_1[i_cpu_address[`INDEX]] <= 0;
          lru_counter_2[i_cpu_address[`INDEX]] <= 1;
          cache_rd_wr_done                     <= 1;
        end
      end
      else
        cache_rd_wr_done <= 0;
    end

    MEM_ACCESS : begin
      cache_rd_wr_done   <= 0;
      if(!valid_1[i_cpu_address[`INDEX]]&i_mem_rd_data_valid&(i_mem_rd_data_tag==i_cpu_address)) begin
        valid_1[i_cpu_address[`INDEX]]  <= 1'b1;
        cache_mem_1[i_cpu_address[`INDEX]] <= i_mem_rd_data;
        dirty_bit_1[i_cpu_address[`INDEX]] <= 1'b0;
        tag_1[i_cpu_address[`INDEX]]       <= i_cpu_address[`TAG];
        //miss                               <= 0;
        mem_rd_wr_done <= 1;
      end
      else if(!valid_2[i_cpu_address[`INDEX]]&i_mem_rd_data_valid&(i_mem_rd_data_tag==i_cpu_address)) begin
        valid_2[i_cpu_address[`INDEX]]  <= 1'b1;
        cache_mem_2[i_cpu_address[`INDEX]] <= i_mem_rd_data;
        dirty_bit_2[i_cpu_address[`INDEX]] <= 1'b0;
        tag_2[i_cpu_address[`INDEX]]       <= i_cpu_address[`TAG];
        //miss                               <= 0;
        mem_rd_wr_done <= 1;
      end
      else if(!lru_counter_1[i_cpu_address[`INDEX]]&i_mem_rd_data_valid&(i_mem_rd_data_tag==i_cpu_address)) begin
        if(dirty_bit_1[i_cpu_address[`INDEX]]) begin
          o_mem_wr_valid  <= 1;
          o_mem_wr_data   <= cache_mem_1[i_cpu_address[`INDEX]];
          o_mem_wr_address <= {tag_1[i_cpu_address[`INDEX]],i_cpu_address[`INDEX],6'd0};          
        end
        cache_mem_1[i_cpu_address[`INDEX]]   <= i_mem_rd_data;
        tag_1[i_cpu_address[`INDEX]]         <= i_cpu_address[`TAG];
        dirty_bit_1[i_cpu_address[`INDEX]]   <= 0;
        //miss <= 0;
        mem_rd_wr_done <= 1;
      end
      else if(!lru_counter_2[i_cpu_address[`INDEX]]&i_mem_rd_data_valid&(i_mem_rd_data_tag==i_cpu_address)) begin
        if(dirty_bit_2[i_cpu_address[`INDEX]]) begin
          o_mem_wr_valid  <= 1;
          o_mem_wr_data   <= cache_mem_2[i_cpu_address[`INDEX]];
          o_mem_wr_address <= {tag_2[i_cpu_address[`INDEX]],i_cpu_address[`INDEX],6'd0};
        end
        cache_mem_2[i_cpu_address[`INDEX]]   <= i_mem_rd_data;
        tag_2[i_cpu_address[`INDEX]]         <= i_cpu_address[`TAG];
        dirty_bit_2[i_cpu_address[`INDEX]]   <= 0;
        //miss <= 0;
        mem_rd_wr_done <= 1;
      end
      else begin
        mem_rd_wr_done <= 0;
      end
    end
    endcase
  end
  else if(~rst_n) begin
    cache_rd_wr_done <=0;
    mem_rd_wr_done   <=0;
    o_cache_busy <=0;
    o_cpu_dout_data <= 0;
    o_cpu_dout_valid <= 0;
    o_mem_wr_address <= 0;
    o_mem_wr_data    <= 0;
    o_mem_wr_valid   <= 0;
    valid_1[0]  <=   0;valid_2[0]  <=   0;dirty_bit_1[0] <= 0;dirty_bit_2[0] <= 0;lru_counter_1[0] <= 0;lru_counter_2[0] <= 0;tag_1[0] <= 0;tag_2[0] <= 0;cache_mem_1[0] <= 0;cache_mem_2[0] <= 0;
    valid_1[1]  <=   0;valid_2[1]  <=   0;dirty_bit_1[1] <= 0;dirty_bit_2[1] <= 0;lru_counter_1[1] <= 0;lru_counter_2[1] <= 0;tag_1[1] <= 0;tag_2[1] <= 0;cache_mem_1[1] <= 0;cache_mem_2[1] <= 0;
    valid_1[2]  <=   0;valid_2[2]  <=   0;dirty_bit_1[2] <= 0;dirty_bit_2[2] <= 0;lru_counter_1[2] <= 0;lru_counter_2[2] <= 0;tag_1[2] <= 0;tag_2[2] <= 0;cache_mem_1[2] <= 0;cache_mem_2[2] <= 0;
    valid_1[3]  <=   0;valid_2[3]  <=   0;dirty_bit_1[3] <= 0;dirty_bit_2[3] <= 0;lru_counter_1[3] <= 0;lru_counter_2[3] <= 0;tag_1[3] <= 0;tag_2[3] <= 0;cache_mem_1[3] <= 0;cache_mem_2[3] <= 0;
    valid_1[4]  <=   0;valid_2[4]  <=   0;dirty_bit_1[4] <= 0;dirty_bit_2[4] <= 0;lru_counter_1[4] <= 0;lru_counter_2[4] <= 0;tag_1[4] <= 0;tag_2[4] <= 0;cache_mem_1[4] <= 0;cache_mem_2[4] <= 0;
    valid_1[5]  <=   0;valid_2[5]  <=   0;dirty_bit_1[5] <= 0;dirty_bit_2[5] <= 0;lru_counter_1[5] <= 0;lru_counter_2[5] <= 0;tag_1[5] <= 0;tag_2[5] <= 0;cache_mem_1[5] <= 0;cache_mem_2[5] <= 0;
    valid_1[6]  <=   0;valid_2[6]  <=   0;dirty_bit_1[6] <= 0;dirty_bit_2[6] <= 0;lru_counter_1[6] <= 0;lru_counter_2[6] <= 0;tag_1[6] <= 0;tag_2[6] <= 0;cache_mem_1[6] <= 0;cache_mem_2[6] <= 0;
    valid_1[7]  <=   0;valid_2[7]  <=   0;dirty_bit_1[7] <= 0;dirty_bit_2[7] <= 0;lru_counter_1[7] <= 0;lru_counter_2[7] <= 0;tag_1[7] <= 0;tag_2[7] <= 0;cache_mem_1[7] <= 0;cache_mem_2[7] <= 0;
    valid_1[8]  <=   0;valid_2[8]  <=   0;dirty_bit_1[8] <= 0;dirty_bit_2[8] <= 0;lru_counter_1[8] <= 0;lru_counter_2[8] <= 0;tag_1[8] <= 0;tag_2[8] <= 0;cache_mem_1[8] <= 0;cache_mem_2[8] <= 0;
    valid_1[9]  <=   0;valid_2[9]  <=   0;dirty_bit_1[9] <= 0;dirty_bit_2[9] <= 0;lru_counter_1[9] <= 0;lru_counter_2[9] <= 0;tag_1[9] <= 0;tag_2[9] <= 0;cache_mem_1[9] <= 0;cache_mem_2[9] <= 0;
    valid_1[10]  <=   0;valid_2[10]  <=   0;dirty_bit_1[10] <= 0;dirty_bit_2[10] <= 0;lru_counter_1[10] <= 0;lru_counter_2[10] <= 0;tag_1[10] <= 0;tag_2[10] <= 0;cache_mem_1[10] <= 0;cache_mem_2[10] <= 0;
    valid_1[11]  <=   0;valid_2[11]  <=   0;dirty_bit_1[11] <= 0;dirty_bit_2[11] <= 0;lru_counter_1[11] <= 0;lru_counter_2[11] <= 0;tag_1[11] <= 0;tag_2[11] <= 0;cache_mem_1[11] <= 0;cache_mem_2[11] <= 0;
    valid_1[12]  <=   0;valid_2[12]  <=   0;dirty_bit_1[12] <= 0;dirty_bit_2[12] <= 0;lru_counter_1[12] <= 0;lru_counter_2[12] <= 0;tag_1[12] <= 0;tag_2[12] <= 0;cache_mem_1[12] <= 0;cache_mem_2[12] <= 0;
    valid_1[13]  <=   0;valid_2[13]  <=   0;dirty_bit_1[13] <= 0;dirty_bit_2[13] <= 0;lru_counter_1[13] <= 0;lru_counter_2[13] <= 0;tag_1[13] <= 0;tag_2[13] <= 0;cache_mem_1[13] <= 0;cache_mem_2[13] <= 0;
    valid_1[14]  <=   0;valid_2[14]  <=   0;dirty_bit_1[14] <= 0;dirty_bit_2[14] <= 0;lru_counter_1[14] <= 0;lru_counter_2[14] <= 0;tag_1[14] <= 0;tag_2[14] <= 0;cache_mem_1[14] <= 0;cache_mem_2[14] <= 0;
    valid_1[15]  <=   0;valid_2[15]  <=   0;dirty_bit_1[15] <= 0;dirty_bit_2[15] <= 0;lru_counter_1[15] <= 0;lru_counter_2[15] <= 0;tag_1[15] <= 0;tag_2[15] <= 0;cache_mem_1[15] <= 0;cache_mem_2[15] <= 0;
    valid_1[16]  <=   0;valid_2[16]  <=   0;dirty_bit_1[16] <= 0;dirty_bit_2[16] <= 0;lru_counter_1[16] <= 0;lru_counter_2[16] <= 0;tag_1[16] <= 0;tag_2[16] <= 0;cache_mem_1[16] <= 0;cache_mem_2[16] <= 0;
    valid_1[17]  <=   0;valid_2[17]  <=   0;dirty_bit_1[17] <= 0;dirty_bit_2[17] <= 0;lru_counter_1[17] <= 0;lru_counter_2[17] <= 0;tag_1[17] <= 0;tag_2[17] <= 0;cache_mem_1[17] <= 0;cache_mem_2[17] <= 0;
    valid_1[18]  <=   0;valid_2[18]  <=   0;dirty_bit_1[18] <= 0;dirty_bit_2[18] <= 0;lru_counter_1[18] <= 0;lru_counter_2[18] <= 0;tag_1[18] <= 0;tag_2[18] <= 0;cache_mem_1[18] <= 0;cache_mem_2[18] <= 0;
    valid_1[19]  <=   0;valid_2[19]  <=   0;dirty_bit_1[19] <= 0;dirty_bit_2[19] <= 0;lru_counter_1[19] <= 0;lru_counter_2[19] <= 0;tag_1[19] <= 0;tag_2[19] <= 0;cache_mem_1[19] <= 0;cache_mem_2[19] <= 0;
    valid_1[20]  <=   0;valid_2[20]  <=   0;dirty_bit_1[20] <= 0;dirty_bit_2[20] <= 0;lru_counter_1[20] <= 0;lru_counter_2[20] <= 0;tag_1[20] <= 0;tag_2[20] <= 0;cache_mem_1[20] <= 0;cache_mem_2[20] <= 0;
    valid_1[21]  <=   0;valid_2[21]  <=   0;dirty_bit_1[21] <= 0;dirty_bit_2[21] <= 0;lru_counter_1[21] <= 0;lru_counter_2[21] <= 0;tag_1[21] <= 0;tag_2[21] <= 0;cache_mem_1[21] <= 0;cache_mem_2[21] <= 0;
    valid_1[22]  <=   0;valid_2[22]  <=   0;dirty_bit_1[22] <= 0;dirty_bit_2[22] <= 0;lru_counter_1[22] <= 0;lru_counter_2[22] <= 0;tag_1[22] <= 0;tag_2[22] <= 0;cache_mem_1[22] <= 0;cache_mem_2[22] <= 0;
    valid_1[23]  <=   0;valid_2[23]  <=   0;dirty_bit_1[23] <= 0;dirty_bit_2[23] <= 0;lru_counter_1[23] <= 0;lru_counter_2[23] <= 0;tag_1[23] <= 0;tag_2[23] <= 0;cache_mem_1[23] <= 0;cache_mem_2[23] <= 0;
    valid_1[24]  <=   0;valid_2[24]  <=   0;dirty_bit_1[24] <= 0;dirty_bit_2[24] <= 0;lru_counter_1[24] <= 0;lru_counter_2[24] <= 0;tag_1[24] <= 0;tag_2[24] <= 0;cache_mem_1[24] <= 0;cache_mem_2[24] <= 0;
    valid_1[25]  <=   0;valid_2[25]  <=   0;dirty_bit_1[25] <= 0;dirty_bit_2[25] <= 0;lru_counter_1[25] <= 0;lru_counter_2[25] <= 0;tag_1[25] <= 0;tag_2[25] <= 0;cache_mem_1[25] <= 0;cache_mem_2[25] <= 0;
    valid_1[26]  <=   0;valid_2[26]  <=   0;dirty_bit_1[26] <= 0;dirty_bit_2[26] <= 0;lru_counter_1[26] <= 0;lru_counter_2[26] <= 0;tag_1[26] <= 0;tag_2[26] <= 0;cache_mem_1[26] <= 0;cache_mem_2[26] <= 0;
    valid_1[27]  <=   0;valid_2[27]  <=   0;dirty_bit_1[27] <= 0;dirty_bit_2[27] <= 0;lru_counter_1[27] <= 0;lru_counter_2[27] <= 0;tag_1[27] <= 0;tag_2[27] <= 0;cache_mem_1[27] <= 0;cache_mem_2[27] <= 0;
    valid_1[28]  <=   0;valid_2[28]  <=   0;dirty_bit_1[28] <= 0;dirty_bit_2[28] <= 0;lru_counter_1[28] <= 0;lru_counter_2[28] <= 0;tag_1[28] <= 0;tag_2[28] <= 0;cache_mem_1[28] <= 0;cache_mem_2[28] <= 0;
    valid_1[29]  <=   0;valid_2[29]  <=   0;dirty_bit_1[29] <= 0;dirty_bit_2[29] <= 0;lru_counter_1[29] <= 0;lru_counter_2[29] <= 0;tag_1[29] <= 0;tag_2[29] <= 0;cache_mem_1[29] <= 0;cache_mem_2[29] <= 0;
    valid_1[30]  <=   0;valid_2[30]  <=   0;dirty_bit_1[30] <= 0;dirty_bit_2[30] <= 0;lru_counter_1[30] <= 0;lru_counter_2[30] <= 0;tag_1[30] <= 0;tag_2[30] <= 0;cache_mem_1[30] <= 0;cache_mem_2[30] <= 0;
    valid_1[31]  <=   0;valid_2[31]  <=   0;dirty_bit_1[31] <= 0;dirty_bit_2[31] <= 0;lru_counter_1[31] <= 0;lru_counter_2[31] <= 0;tag_1[31] <= 0;tag_2[31] <= 0;cache_mem_1[31] <= 0;cache_mem_2[31] <= 0;
    valid_1[32]  <=   0;valid_2[32]  <=   0;dirty_bit_1[32] <= 0;dirty_bit_2[32] <= 0;lru_counter_1[32] <= 0;lru_counter_2[32] <= 0;tag_1[32] <= 0;tag_2[32] <= 0;cache_mem_1[32] <= 0;cache_mem_2[32] <= 0;
    valid_1[33]  <=   0;valid_2[33]  <=   0;dirty_bit_1[33] <= 0;dirty_bit_2[33] <= 0;lru_counter_1[33] <= 0;lru_counter_2[33] <= 0;tag_1[33] <= 0;tag_2[33] <= 0;cache_mem_1[33] <= 0;cache_mem_2[33] <= 0;
    valid_1[34]  <=   0;valid_2[34]  <=   0;dirty_bit_1[34] <= 0;dirty_bit_2[34] <= 0;lru_counter_1[34] <= 0;lru_counter_2[34] <= 0;tag_1[34] <= 0;tag_2[34] <= 0;cache_mem_1[34] <= 0;cache_mem_2[34] <= 0;
    valid_1[35]  <=   0;valid_2[35]  <=   0;dirty_bit_1[35] <= 0;dirty_bit_2[35] <= 0;lru_counter_1[35] <= 0;lru_counter_2[35] <= 0;tag_1[35] <= 0;tag_2[35] <= 0;cache_mem_1[35] <= 0;cache_mem_2[35] <= 0;
    valid_1[36]  <=   0;valid_2[36]  <=   0;dirty_bit_1[36] <= 0;dirty_bit_2[36] <= 0;lru_counter_1[36] <= 0;lru_counter_2[36] <= 0;tag_1[36] <= 0;tag_2[36] <= 0;cache_mem_1[36] <= 0;cache_mem_2[36] <= 0;
    valid_1[37]  <=   0;valid_2[37]  <=   0;dirty_bit_1[37] <= 0;dirty_bit_2[37] <= 0;lru_counter_1[37] <= 0;lru_counter_2[37] <= 0;tag_1[37] <= 0;tag_2[37] <= 0;cache_mem_1[37] <= 0;cache_mem_2[37] <= 0;
    valid_1[38]  <=   0;valid_2[38]  <=   0;dirty_bit_1[38] <= 0;dirty_bit_2[38] <= 0;lru_counter_1[38] <= 0;lru_counter_2[38] <= 0;tag_1[38] <= 0;tag_2[38] <= 0;cache_mem_1[38] <= 0;cache_mem_2[38] <= 0;
    valid_1[39]  <=   0;valid_2[39]  <=   0;dirty_bit_1[39] <= 0;dirty_bit_2[39] <= 0;lru_counter_1[39] <= 0;lru_counter_2[39] <= 0;tag_1[39] <= 0;tag_2[39] <= 0;cache_mem_1[39] <= 0;cache_mem_2[39] <= 0;
    valid_1[40]  <=   0;valid_2[40]  <=   0;dirty_bit_1[40] <= 0;dirty_bit_2[40] <= 0;lru_counter_1[40] <= 0;lru_counter_2[40] <= 0;tag_1[40] <= 0;tag_2[40] <= 0;cache_mem_1[40] <= 0;cache_mem_2[40] <= 0;
    valid_1[41]  <=   0;valid_2[41]  <=   0;dirty_bit_1[41] <= 0;dirty_bit_2[41] <= 0;lru_counter_1[41] <= 0;lru_counter_2[41] <= 0;tag_1[41] <= 0;tag_2[41] <= 0;cache_mem_1[41] <= 0;cache_mem_2[41] <= 0;
    valid_1[42]  <=   0;valid_2[42]  <=   0;dirty_bit_1[42] <= 0;dirty_bit_2[42] <= 0;lru_counter_1[42] <= 0;lru_counter_2[42] <= 0;tag_1[42] <= 0;tag_2[42] <= 0;cache_mem_1[42] <= 0;cache_mem_2[42] <= 0;
    valid_1[43]  <=   0;valid_2[43]  <=   0;dirty_bit_1[43] <= 0;dirty_bit_2[43] <= 0;lru_counter_1[43] <= 0;lru_counter_2[43] <= 0;tag_1[43] <= 0;tag_2[43] <= 0;cache_mem_1[43] <= 0;cache_mem_2[43] <= 0;
    valid_1[44]  <=   0;valid_2[44]  <=   0;dirty_bit_1[44] <= 0;dirty_bit_2[44] <= 0;lru_counter_1[44] <= 0;lru_counter_2[44] <= 0;tag_1[44] <= 0;tag_2[44] <= 0;cache_mem_1[44] <= 0;cache_mem_2[44] <= 0;
    valid_1[45]  <=   0;valid_2[45]  <=   0;dirty_bit_1[45] <= 0;dirty_bit_2[45] <= 0;lru_counter_1[45] <= 0;lru_counter_2[45] <= 0;tag_1[45] <= 0;tag_2[45] <= 0;cache_mem_1[45] <= 0;cache_mem_2[45] <= 0;
    valid_1[46]  <=   0;valid_2[46]  <=   0;dirty_bit_1[46] <= 0;dirty_bit_2[46] <= 0;lru_counter_1[46] <= 0;lru_counter_2[46] <= 0;tag_1[46] <= 0;tag_2[46] <= 0;cache_mem_1[46] <= 0;cache_mem_2[46] <= 0;
    valid_1[47]  <=   0;valid_2[47]  <=   0;dirty_bit_1[47] <= 0;dirty_bit_2[47] <= 0;lru_counter_1[47] <= 0;lru_counter_2[47] <= 0;tag_1[47] <= 0;tag_2[47] <= 0;cache_mem_1[47] <= 0;cache_mem_2[47] <= 0;
    valid_1[48]  <=   0;valid_2[48]  <=   0;dirty_bit_1[48] <= 0;dirty_bit_2[48] <= 0;lru_counter_1[48] <= 0;lru_counter_2[48] <= 0;tag_1[48] <= 0;tag_2[48] <= 0;cache_mem_1[48] <= 0;cache_mem_2[48] <= 0;
    valid_1[49]  <=   0;valid_2[49]  <=   0;dirty_bit_1[49] <= 0;dirty_bit_2[49] <= 0;lru_counter_1[49] <= 0;lru_counter_2[49] <= 0;tag_1[49] <= 0;tag_2[49] <= 0;cache_mem_1[49] <= 0;cache_mem_2[49] <= 0;
    valid_1[50]  <=   0;valid_2[50]  <=   0;dirty_bit_1[50] <= 0;dirty_bit_2[50] <= 0;lru_counter_1[50] <= 0;lru_counter_2[50] <= 0;tag_1[50] <= 0;tag_2[50] <= 0;cache_mem_1[50] <= 0;cache_mem_2[50] <= 0;
    valid_1[51]  <=   0;valid_2[51]  <=   0;dirty_bit_1[51] <= 0;dirty_bit_2[51] <= 0;lru_counter_1[51] <= 0;lru_counter_2[51] <= 0;tag_1[51] <= 0;tag_2[51] <= 0;cache_mem_1[51] <= 0;cache_mem_2[51] <= 0;
    valid_1[52]  <=   0;valid_2[52]  <=   0;dirty_bit_1[52] <= 0;dirty_bit_2[52] <= 0;lru_counter_1[52] <= 0;lru_counter_2[52] <= 0;tag_1[52] <= 0;tag_2[52] <= 0;cache_mem_1[52] <= 0;cache_mem_2[52] <= 0;
    valid_1[53]  <=   0;valid_2[53]  <=   0;dirty_bit_1[53] <= 0;dirty_bit_2[53] <= 0;lru_counter_1[53] <= 0;lru_counter_2[53] <= 0;tag_1[53] <= 0;tag_2[53] <= 0;cache_mem_1[53] <= 0;cache_mem_2[53] <= 0;
    valid_1[54]  <=   0;valid_2[54]  <=   0;dirty_bit_1[54] <= 0;dirty_bit_2[54] <= 0;lru_counter_1[54] <= 0;lru_counter_2[54] <= 0;tag_1[54] <= 0;tag_2[54] <= 0;cache_mem_1[54] <= 0;cache_mem_2[54] <= 0;
    valid_1[55]  <=   0;valid_2[55]  <=   0;dirty_bit_1[55] <= 0;dirty_bit_2[55] <= 0;lru_counter_1[55] <= 0;lru_counter_2[55] <= 0;tag_1[55] <= 0;tag_2[55] <= 0;cache_mem_1[55] <= 0;cache_mem_2[55] <= 0;
    valid_1[56]  <=   0;valid_2[56]  <=   0;dirty_bit_1[56] <= 0;dirty_bit_2[56] <= 0;lru_counter_1[56] <= 0;lru_counter_2[56] <= 0;tag_1[56] <= 0;tag_2[56] <= 0;cache_mem_1[56] <= 0;cache_mem_2[56] <= 0;
    valid_1[57]  <=   0;valid_2[57]  <=   0;dirty_bit_1[57] <= 0;dirty_bit_2[57] <= 0;lru_counter_1[57] <= 0;lru_counter_2[57] <= 0;tag_1[57] <= 0;tag_2[57] <= 0;cache_mem_1[57] <= 0;cache_mem_2[57] <= 0;
    valid_1[58]  <=   0;valid_2[58]  <=   0;dirty_bit_1[58] <= 0;dirty_bit_2[58] <= 0;lru_counter_1[58] <= 0;lru_counter_2[58] <= 0;tag_1[58] <= 0;tag_2[58] <= 0;cache_mem_1[58] <= 0;cache_mem_2[58] <= 0;
    valid_1[59]  <=   0;valid_2[59]  <=   0;dirty_bit_1[59] <= 0;dirty_bit_2[59] <= 0;lru_counter_1[59] <= 0;lru_counter_2[59] <= 0;tag_1[59] <= 0;tag_2[59] <= 0;cache_mem_1[59] <= 0;cache_mem_2[59] <= 0;
    valid_1[60]  <=   0;valid_2[60]  <=   0;dirty_bit_1[60] <= 0;dirty_bit_2[60] <= 0;lru_counter_1[60] <= 0;lru_counter_2[60] <= 0;tag_1[60] <= 0;tag_2[60] <= 0;cache_mem_1[60] <= 0;cache_mem_2[60] <= 0;
    valid_1[61]  <=   0;valid_2[61]  <=   0;dirty_bit_1[61] <= 0;dirty_bit_2[61] <= 0;lru_counter_1[61] <= 0;lru_counter_2[61] <= 0;tag_1[61] <= 0;tag_2[61] <= 0;cache_mem_1[61] <= 0;cache_mem_2[61] <= 0;
    valid_1[62]  <=   0;valid_2[62]  <=   0;dirty_bit_1[62] <= 0;dirty_bit_2[62] <= 0;lru_counter_1[62] <= 0;lru_counter_2[62] <= 0;tag_1[62] <= 0;tag_2[62] <= 0;cache_mem_1[62] <= 0;cache_mem_2[62] <= 0;
    valid_1[63]  <=   0;valid_2[63]  <=   0;dirty_bit_1[63] <= 0;dirty_bit_2[63] <= 0;lru_counter_1[63] <= 0;lru_counter_2[63] <= 0;tag_1[63] <= 0;tag_2[63] <= 0;cache_mem_1[63] <= 0;cache_mem_2[63] <= 0;
    valid_1[64]  <=   0;valid_2[64]  <=   0;dirty_bit_1[64] <= 0;dirty_bit_2[64] <= 0;lru_counter_1[64] <= 0;lru_counter_2[64] <= 0;tag_1[64] <= 0;tag_2[64] <= 0;cache_mem_1[64] <= 0;cache_mem_2[64] <= 0;
    valid_1[65]  <=   0;valid_2[65]  <=   0;dirty_bit_1[65] <= 0;dirty_bit_2[65] <= 0;lru_counter_1[65] <= 0;lru_counter_2[65] <= 0;tag_1[65] <= 0;tag_2[65] <= 0;cache_mem_1[65] <= 0;cache_mem_2[65] <= 0;
    valid_1[66]  <=   0;valid_2[66]  <=   0;dirty_bit_1[66] <= 0;dirty_bit_2[66] <= 0;lru_counter_1[66] <= 0;lru_counter_2[66] <= 0;tag_1[66] <= 0;tag_2[66] <= 0;cache_mem_1[66] <= 0;cache_mem_2[66] <= 0;
    valid_1[67]  <=   0;valid_2[67]  <=   0;dirty_bit_1[67] <= 0;dirty_bit_2[67] <= 0;lru_counter_1[67] <= 0;lru_counter_2[67] <= 0;tag_1[67] <= 0;tag_2[67] <= 0;cache_mem_1[67] <= 0;cache_mem_2[67] <= 0;
    valid_1[68]  <=   0;valid_2[68]  <=   0;dirty_bit_1[68] <= 0;dirty_bit_2[68] <= 0;lru_counter_1[68] <= 0;lru_counter_2[68] <= 0;tag_1[68] <= 0;tag_2[68] <= 0;cache_mem_1[68] <= 0;cache_mem_2[68] <= 0;
    valid_1[69]  <=   0;valid_2[69]  <=   0;dirty_bit_1[69] <= 0;dirty_bit_2[69] <= 0;lru_counter_1[69] <= 0;lru_counter_2[69] <= 0;tag_1[69] <= 0;tag_2[69] <= 0;cache_mem_1[69] <= 0;cache_mem_2[69] <= 0;
    valid_1[70]  <=   0;valid_2[70]  <=   0;dirty_bit_1[70] <= 0;dirty_bit_2[70] <= 0;lru_counter_1[70] <= 0;lru_counter_2[70] <= 0;tag_1[70] <= 0;tag_2[70] <= 0;cache_mem_1[70] <= 0;cache_mem_2[70] <= 0;
    valid_1[71]  <=   0;valid_2[71]  <=   0;dirty_bit_1[71] <= 0;dirty_bit_2[71] <= 0;lru_counter_1[71] <= 0;lru_counter_2[71] <= 0;tag_1[71] <= 0;tag_2[71] <= 0;cache_mem_1[71] <= 0;cache_mem_2[71] <= 0;
    valid_1[72]  <=   0;valid_2[72]  <=   0;dirty_bit_1[72] <= 0;dirty_bit_2[72] <= 0;lru_counter_1[72] <= 0;lru_counter_2[72] <= 0;tag_1[72] <= 0;tag_2[72] <= 0;cache_mem_1[72] <= 0;cache_mem_2[72] <= 0;
    valid_1[73]  <=   0;valid_2[73]  <=   0;dirty_bit_1[73] <= 0;dirty_bit_2[73] <= 0;lru_counter_1[73] <= 0;lru_counter_2[73] <= 0;tag_1[73] <= 0;tag_2[73] <= 0;cache_mem_1[73] <= 0;cache_mem_2[73] <= 0;
    valid_1[74]  <=   0;valid_2[74]  <=   0;dirty_bit_1[74] <= 0;dirty_bit_2[74] <= 0;lru_counter_1[74] <= 0;lru_counter_2[74] <= 0;tag_1[74] <= 0;tag_2[74] <= 0;cache_mem_1[74] <= 0;cache_mem_2[74] <= 0;
    valid_1[75]  <=   0;valid_2[75]  <=   0;dirty_bit_1[75] <= 0;dirty_bit_2[75] <= 0;lru_counter_1[75] <= 0;lru_counter_2[75] <= 0;tag_1[75] <= 0;tag_2[75] <= 0;cache_mem_1[75] <= 0;cache_mem_2[75] <= 0;
    valid_1[76]  <=   0;valid_2[76]  <=   0;dirty_bit_1[76] <= 0;dirty_bit_2[76] <= 0;lru_counter_1[76] <= 0;lru_counter_2[76] <= 0;tag_1[76] <= 0;tag_2[76] <= 0;cache_mem_1[76] <= 0;cache_mem_2[76] <= 0;
    valid_1[77]  <=   0;valid_2[77]  <=   0;dirty_bit_1[77] <= 0;dirty_bit_2[77] <= 0;lru_counter_1[77] <= 0;lru_counter_2[77] <= 0;tag_1[77] <= 0;tag_2[77] <= 0;cache_mem_1[77] <= 0;cache_mem_2[77] <= 0;
    valid_1[78]  <=   0;valid_2[78]  <=   0;dirty_bit_1[78] <= 0;dirty_bit_2[78] <= 0;lru_counter_1[78] <= 0;lru_counter_2[78] <= 0;tag_1[78] <= 0;tag_2[78] <= 0;cache_mem_1[78] <= 0;cache_mem_2[78] <= 0;
    valid_1[79]  <=   0;valid_2[79]  <=   0;dirty_bit_1[79] <= 0;dirty_bit_2[79] <= 0;lru_counter_1[79] <= 0;lru_counter_2[79] <= 0;tag_1[79] <= 0;tag_2[79] <= 0;cache_mem_1[79] <= 0;cache_mem_2[79] <= 0;
    valid_1[80]  <=   0;valid_2[80]  <=   0;dirty_bit_1[80] <= 0;dirty_bit_2[80] <= 0;lru_counter_1[80] <= 0;lru_counter_2[80] <= 0;tag_1[80] <= 0;tag_2[80] <= 0;cache_mem_1[80] <= 0;cache_mem_2[80] <= 0;
    valid_1[81]  <=   0;valid_2[81]  <=   0;dirty_bit_1[81] <= 0;dirty_bit_2[81] <= 0;lru_counter_1[81] <= 0;lru_counter_2[81] <= 0;tag_1[81] <= 0;tag_2[81] <= 0;cache_mem_1[81] <= 0;cache_mem_2[81] <= 0;
    valid_1[82]  <=   0;valid_2[82]  <=   0;dirty_bit_1[82] <= 0;dirty_bit_2[82] <= 0;lru_counter_1[82] <= 0;lru_counter_2[82] <= 0;tag_1[82] <= 0;tag_2[82] <= 0;cache_mem_1[82] <= 0;cache_mem_2[82] <= 0;
    valid_1[83]  <=   0;valid_2[83]  <=   0;dirty_bit_1[83] <= 0;dirty_bit_2[83] <= 0;lru_counter_1[83] <= 0;lru_counter_2[83] <= 0;tag_1[83] <= 0;tag_2[83] <= 0;cache_mem_1[83] <= 0;cache_mem_2[83] <= 0;
    valid_1[84]  <=   0;valid_2[84]  <=   0;dirty_bit_1[84] <= 0;dirty_bit_2[84] <= 0;lru_counter_1[84] <= 0;lru_counter_2[84] <= 0;tag_1[84] <= 0;tag_2[84] <= 0;cache_mem_1[84] <= 0;cache_mem_2[84] <= 0;
    valid_1[85]  <=   0;valid_2[85]  <=   0;dirty_bit_1[85] <= 0;dirty_bit_2[85] <= 0;lru_counter_1[85] <= 0;lru_counter_2[85] <= 0;tag_1[85] <= 0;tag_2[85] <= 0;cache_mem_1[85] <= 0;cache_mem_2[85] <= 0;
    valid_1[86]  <=   0;valid_2[86]  <=   0;dirty_bit_1[86] <= 0;dirty_bit_2[86] <= 0;lru_counter_1[86] <= 0;lru_counter_2[86] <= 0;tag_1[86] <= 0;tag_2[86] <= 0;cache_mem_1[86] <= 0;cache_mem_2[86] <= 0;
    valid_1[87]  <=   0;valid_2[87]  <=   0;dirty_bit_1[87] <= 0;dirty_bit_2[87] <= 0;lru_counter_1[87] <= 0;lru_counter_2[87] <= 0;tag_1[87] <= 0;tag_2[87] <= 0;cache_mem_1[87] <= 0;cache_mem_2[87] <= 0;
    valid_1[88]  <=   0;valid_2[88]  <=   0;dirty_bit_1[88] <= 0;dirty_bit_2[88] <= 0;lru_counter_1[88] <= 0;lru_counter_2[88] <= 0;tag_1[88] <= 0;tag_2[88] <= 0;cache_mem_1[88] <= 0;cache_mem_2[88] <= 0;
    valid_1[89]  <=   0;valid_2[89]  <=   0;dirty_bit_1[89] <= 0;dirty_bit_2[89] <= 0;lru_counter_1[89] <= 0;lru_counter_2[89] <= 0;tag_1[89] <= 0;tag_2[89] <= 0;cache_mem_1[89] <= 0;cache_mem_2[89] <= 0;
    valid_1[90]  <=   0;valid_2[90]  <=   0;dirty_bit_1[90] <= 0;dirty_bit_2[90] <= 0;lru_counter_1[90] <= 0;lru_counter_2[90] <= 0;tag_1[90] <= 0;tag_2[90] <= 0;cache_mem_1[90] <= 0;cache_mem_2[90] <= 0;
    valid_1[91]  <=   0;valid_2[91]  <=   0;dirty_bit_1[91] <= 0;dirty_bit_2[91] <= 0;lru_counter_1[91] <= 0;lru_counter_2[91] <= 0;tag_1[91] <= 0;tag_2[91] <= 0;cache_mem_1[91] <= 0;cache_mem_2[91] <= 0;
    valid_1[92]  <=   0;valid_2[92]  <=   0;dirty_bit_1[92] <= 0;dirty_bit_2[92] <= 0;lru_counter_1[92] <= 0;lru_counter_2[92] <= 0;tag_1[92] <= 0;tag_2[92] <= 0;cache_mem_1[92] <= 0;cache_mem_2[92] <= 0;
    valid_1[93]  <=   0;valid_2[93]  <=   0;dirty_bit_1[93] <= 0;dirty_bit_2[93] <= 0;lru_counter_1[93] <= 0;lru_counter_2[93] <= 0;tag_1[93] <= 0;tag_2[93] <= 0;cache_mem_1[93] <= 0;cache_mem_2[93] <= 0;
    valid_1[94]  <=   0;valid_2[94]  <=   0;dirty_bit_1[94] <= 0;dirty_bit_2[94] <= 0;lru_counter_1[94] <= 0;lru_counter_2[94] <= 0;tag_1[94] <= 0;tag_2[94] <= 0;cache_mem_1[94] <= 0;cache_mem_2[94] <= 0;
    valid_1[95]  <=   0;valid_2[95]  <=   0;dirty_bit_1[95] <= 0;dirty_bit_2[95] <= 0;lru_counter_1[95] <= 0;lru_counter_2[95] <= 0;tag_1[95] <= 0;tag_2[95] <= 0;cache_mem_1[95] <= 0;cache_mem_2[95] <= 0;
    valid_1[96]  <=   0;valid_2[96]  <=   0;dirty_bit_1[96] <= 0;dirty_bit_2[96] <= 0;lru_counter_1[96] <= 0;lru_counter_2[96] <= 0;tag_1[96] <= 0;tag_2[96] <= 0;cache_mem_1[96] <= 0;cache_mem_2[96] <= 0;
    valid_1[97]  <=   0;valid_2[97]  <=   0;dirty_bit_1[97] <= 0;dirty_bit_2[97] <= 0;lru_counter_1[97] <= 0;lru_counter_2[97] <= 0;tag_1[97] <= 0;tag_2[97] <= 0;cache_mem_1[97] <= 0;cache_mem_2[97] <= 0;
    valid_1[98]  <=   0;valid_2[98]  <=   0;dirty_bit_1[98] <= 0;dirty_bit_2[98] <= 0;lru_counter_1[98] <= 0;lru_counter_2[98] <= 0;tag_1[98] <= 0;tag_2[98] <= 0;cache_mem_1[98] <= 0;cache_mem_2[98] <= 0;
    valid_1[99]  <=   0;valid_2[99]  <=   0;dirty_bit_1[99] <= 0;dirty_bit_2[99] <= 0;lru_counter_1[99] <= 0;lru_counter_2[99] <= 0;tag_1[99] <= 0;tag_2[99] <= 0;cache_mem_1[99] <= 0;cache_mem_2[99] <= 0;
    valid_1[100]  <=   0;valid_2[100]  <=   0;dirty_bit_1[100] <= 0;dirty_bit_2[100] <= 0;lru_counter_1[100] <= 0;lru_counter_2[100] <= 0;tag_1[100] <= 0;tag_2[100] <= 0;cache_mem_1[100] <= 0;cache_mem_2[100] <= 0;
    valid_1[101]  <=   0;valid_2[101]  <=   0;dirty_bit_1[101] <= 0;dirty_bit_2[101] <= 0;lru_counter_1[101] <= 0;lru_counter_2[101] <= 0;tag_1[101] <= 0;tag_2[101] <= 0;cache_mem_1[101] <= 0;cache_mem_2[101] <= 0;
    valid_1[102]  <=   0;valid_2[102]  <=   0;dirty_bit_1[102] <= 0;dirty_bit_2[102] <= 0;lru_counter_1[102] <= 0;lru_counter_2[102] <= 0;tag_1[102] <= 0;tag_2[102] <= 0;cache_mem_1[102] <= 0;cache_mem_2[102] <= 0;
    valid_1[103]  <=   0;valid_2[103]  <=   0;dirty_bit_1[103] <= 0;dirty_bit_2[103] <= 0;lru_counter_1[103] <= 0;lru_counter_2[103] <= 0;tag_1[103] <= 0;tag_2[103] <= 0;cache_mem_1[103] <= 0;cache_mem_2[103] <= 0;
    valid_1[104]  <=   0;valid_2[104]  <=   0;dirty_bit_1[104] <= 0;dirty_bit_2[104] <= 0;lru_counter_1[104] <= 0;lru_counter_2[104] <= 0;tag_1[104] <= 0;tag_2[104] <= 0;cache_mem_1[104] <= 0;cache_mem_2[104] <= 0;
    valid_1[105]  <=   0;valid_2[105]  <=   0;dirty_bit_1[105] <= 0;dirty_bit_2[105] <= 0;lru_counter_1[105] <= 0;lru_counter_2[105] <= 0;tag_1[105] <= 0;tag_2[105] <= 0;cache_mem_1[105] <= 0;cache_mem_2[105] <= 0;
    valid_1[106]  <=   0;valid_2[106]  <=   0;dirty_bit_1[106] <= 0;dirty_bit_2[106] <= 0;lru_counter_1[106] <= 0;lru_counter_2[106] <= 0;tag_1[106] <= 0;tag_2[106] <= 0;cache_mem_1[106] <= 0;cache_mem_2[106] <= 0;
    valid_1[107]  <=   0;valid_2[107]  <=   0;dirty_bit_1[107] <= 0;dirty_bit_2[107] <= 0;lru_counter_1[107] <= 0;lru_counter_2[107] <= 0;tag_1[107] <= 0;tag_2[107] <= 0;cache_mem_1[107] <= 0;cache_mem_2[107] <= 0;
    valid_1[108]  <=   0;valid_2[108]  <=   0;dirty_bit_1[108] <= 0;dirty_bit_2[108] <= 0;lru_counter_1[108] <= 0;lru_counter_2[108] <= 0;tag_1[108] <= 0;tag_2[108] <= 0;cache_mem_1[108] <= 0;cache_mem_2[108] <= 0;
    valid_1[109]  <=   0;valid_2[109]  <=   0;dirty_bit_1[109] <= 0;dirty_bit_2[109] <= 0;lru_counter_1[109] <= 0;lru_counter_2[109] <= 0;tag_1[109] <= 0;tag_2[109] <= 0;cache_mem_1[109] <= 0;cache_mem_2[109] <= 0;
    valid_1[110]  <=   0;valid_2[110]  <=   0;dirty_bit_1[110] <= 0;dirty_bit_2[110] <= 0;lru_counter_1[110] <= 0;lru_counter_2[110] <= 0;tag_1[110] <= 0;tag_2[110] <= 0;cache_mem_1[110] <= 0;cache_mem_2[110] <= 0;
    valid_1[111]  <=   0;valid_2[111]  <=   0;dirty_bit_1[111] <= 0;dirty_bit_2[111] <= 0;lru_counter_1[111] <= 0;lru_counter_2[111] <= 0;tag_1[111] <= 0;tag_2[111] <= 0;cache_mem_1[111] <= 0;cache_mem_2[111] <= 0;
    valid_1[112]  <=   0;valid_2[112]  <=   0;dirty_bit_1[112] <= 0;dirty_bit_2[112] <= 0;lru_counter_1[112] <= 0;lru_counter_2[112] <= 0;tag_1[112] <= 0;tag_2[112] <= 0;cache_mem_1[112] <= 0;cache_mem_2[112] <= 0;
    valid_1[113]  <=   0;valid_2[113]  <=   0;dirty_bit_1[113] <= 0;dirty_bit_2[113] <= 0;lru_counter_1[113] <= 0;lru_counter_2[113] <= 0;tag_1[113] <= 0;tag_2[113] <= 0;cache_mem_1[113] <= 0;cache_mem_2[113] <= 0;
    valid_1[114]  <=   0;valid_2[114]  <=   0;dirty_bit_1[114] <= 0;dirty_bit_2[114] <= 0;lru_counter_1[114] <= 0;lru_counter_2[114] <= 0;tag_1[114] <= 0;tag_2[114] <= 0;cache_mem_1[114] <= 0;cache_mem_2[114] <= 0;
    valid_1[115]  <=   0;valid_2[115]  <=   0;dirty_bit_1[115] <= 0;dirty_bit_2[115] <= 0;lru_counter_1[115] <= 0;lru_counter_2[115] <= 0;tag_1[115] <= 0;tag_2[115] <= 0;cache_mem_1[115] <= 0;cache_mem_2[115] <= 0;
    valid_1[116]  <=   0;valid_2[116]  <=   0;dirty_bit_1[116] <= 0;dirty_bit_2[116] <= 0;lru_counter_1[116] <= 0;lru_counter_2[116] <= 0;tag_1[116] <= 0;tag_2[116] <= 0;cache_mem_1[116] <= 0;cache_mem_2[116] <= 0;
    valid_1[117]  <=   0;valid_2[117]  <=   0;dirty_bit_1[117] <= 0;dirty_bit_2[117] <= 0;lru_counter_1[117] <= 0;lru_counter_2[117] <= 0;tag_1[117] <= 0;tag_2[117] <= 0;cache_mem_1[117] <= 0;cache_mem_2[117] <= 0;
    valid_1[118]  <=   0;valid_2[118]  <=   0;dirty_bit_1[118] <= 0;dirty_bit_2[118] <= 0;lru_counter_1[118] <= 0;lru_counter_2[118] <= 0;tag_1[118] <= 0;tag_2[118] <= 0;cache_mem_1[118] <= 0;cache_mem_2[118] <= 0;
    valid_1[119]  <=   0;valid_2[119]  <=   0;dirty_bit_1[119] <= 0;dirty_bit_2[119] <= 0;lru_counter_1[119] <= 0;lru_counter_2[119] <= 0;tag_1[119] <= 0;tag_2[119] <= 0;cache_mem_1[119] <= 0;cache_mem_2[119] <= 0;
    valid_1[120]  <=   0;valid_2[120]  <=   0;dirty_bit_1[120] <= 0;dirty_bit_2[120] <= 0;lru_counter_1[120] <= 0;lru_counter_2[120] <= 0;tag_1[120] <= 0;tag_2[120] <= 0;cache_mem_1[120] <= 0;cache_mem_2[120] <= 0;
    valid_1[121]  <=   0;valid_2[121]  <=   0;dirty_bit_1[121] <= 0;dirty_bit_2[121] <= 0;lru_counter_1[121] <= 0;lru_counter_2[121] <= 0;tag_1[121] <= 0;tag_2[121] <= 0;cache_mem_1[121] <= 0;cache_mem_2[121] <= 0;
    valid_1[122]  <=   0;valid_2[122]  <=   0;dirty_bit_1[122] <= 0;dirty_bit_2[122] <= 0;lru_counter_1[122] <= 0;lru_counter_2[122] <= 0;tag_1[122] <= 0;tag_2[122] <= 0;cache_mem_1[122] <= 0;cache_mem_2[122] <= 0;
    valid_1[123]  <=   0;valid_2[123]  <=   0;dirty_bit_1[123] <= 0;dirty_bit_2[123] <= 0;lru_counter_1[123] <= 0;lru_counter_2[123] <= 0;tag_1[123] <= 0;tag_2[123] <= 0;cache_mem_1[123] <= 0;cache_mem_2[123] <= 0;
    valid_1[124]  <=   0;valid_2[124]  <=   0;dirty_bit_1[124] <= 0;dirty_bit_2[124] <= 0;lru_counter_1[124] <= 0;lru_counter_2[124] <= 0;tag_1[124] <= 0;tag_2[124] <= 0;cache_mem_1[124] <= 0;cache_mem_2[124] <= 0;
    valid_1[125]  <=   0;valid_2[125]  <=   0;dirty_bit_1[125] <= 0;dirty_bit_2[125] <= 0;lru_counter_1[125] <= 0;lru_counter_2[125] <= 0;tag_1[125] <= 0;tag_2[125] <= 0;cache_mem_1[125] <= 0;cache_mem_2[125] <= 0;
    valid_1[126]  <=   0;valid_2[126]  <=   0;dirty_bit_1[126] <= 0;dirty_bit_2[126] <= 0;lru_counter_1[126] <= 0;lru_counter_2[126] <= 0;tag_1[126] <= 0;tag_2[126] <= 0;cache_mem_1[126] <= 0;cache_mem_2[126] <= 0;
    valid_1[127]  <=   0;valid_2[127]  <=   0;dirty_bit_1[127] <= 0;dirty_bit_2[127] <= 0;lru_counter_1[127] <= 0;lru_counter_2[127] <= 0;tag_1[127] <= 0;tag_2[127] <= 0;cache_mem_1[127] <= 0;cache_mem_2[127] <= 0;
    valid_1[128]  <=   0;valid_2[128]  <=   0;dirty_bit_1[128] <= 0;dirty_bit_2[128] <= 0;lru_counter_1[128] <= 0;lru_counter_2[128] <= 0;tag_1[128] <= 0;tag_2[128] <= 0;cache_mem_1[128] <= 0;cache_mem_2[128] <= 0;
    valid_1[129]  <=   0;valid_2[129]  <=   0;dirty_bit_1[129] <= 0;dirty_bit_2[129] <= 0;lru_counter_1[129] <= 0;lru_counter_2[129] <= 0;tag_1[129] <= 0;tag_2[129] <= 0;cache_mem_1[129] <= 0;cache_mem_2[129] <= 0;
    valid_1[130]  <=   0;valid_2[130]  <=   0;dirty_bit_1[130] <= 0;dirty_bit_2[130] <= 0;lru_counter_1[130] <= 0;lru_counter_2[130] <= 0;tag_1[130] <= 0;tag_2[130] <= 0;cache_mem_1[130] <= 0;cache_mem_2[130] <= 0;
    valid_1[131]  <=   0;valid_2[131]  <=   0;dirty_bit_1[131] <= 0;dirty_bit_2[131] <= 0;lru_counter_1[131] <= 0;lru_counter_2[131] <= 0;tag_1[131] <= 0;tag_2[131] <= 0;cache_mem_1[131] <= 0;cache_mem_2[131] <= 0;
    valid_1[132]  <=   0;valid_2[132]  <=   0;dirty_bit_1[132] <= 0;dirty_bit_2[132] <= 0;lru_counter_1[132] <= 0;lru_counter_2[132] <= 0;tag_1[132] <= 0;tag_2[132] <= 0;cache_mem_1[132] <= 0;cache_mem_2[132] <= 0;
    valid_1[133]  <=   0;valid_2[133]  <=   0;dirty_bit_1[133] <= 0;dirty_bit_2[133] <= 0;lru_counter_1[133] <= 0;lru_counter_2[133] <= 0;tag_1[133] <= 0;tag_2[133] <= 0;cache_mem_1[133] <= 0;cache_mem_2[133] <= 0;
    valid_1[134]  <=   0;valid_2[134]  <=   0;dirty_bit_1[134] <= 0;dirty_bit_2[134] <= 0;lru_counter_1[134] <= 0;lru_counter_2[134] <= 0;tag_1[134] <= 0;tag_2[134] <= 0;cache_mem_1[134] <= 0;cache_mem_2[134] <= 0;
    valid_1[135]  <=   0;valid_2[135]  <=   0;dirty_bit_1[135] <= 0;dirty_bit_2[135] <= 0;lru_counter_1[135] <= 0;lru_counter_2[135] <= 0;tag_1[135] <= 0;tag_2[135] <= 0;cache_mem_1[135] <= 0;cache_mem_2[135] <= 0;
    valid_1[136]  <=   0;valid_2[136]  <=   0;dirty_bit_1[136] <= 0;dirty_bit_2[136] <= 0;lru_counter_1[136] <= 0;lru_counter_2[136] <= 0;tag_1[136] <= 0;tag_2[136] <= 0;cache_mem_1[136] <= 0;cache_mem_2[136] <= 0;
    valid_1[137]  <=   0;valid_2[137]  <=   0;dirty_bit_1[137] <= 0;dirty_bit_2[137] <= 0;lru_counter_1[137] <= 0;lru_counter_2[137] <= 0;tag_1[137] <= 0;tag_2[137] <= 0;cache_mem_1[137] <= 0;cache_mem_2[137] <= 0;
    valid_1[138]  <=   0;valid_2[138]  <=   0;dirty_bit_1[138] <= 0;dirty_bit_2[138] <= 0;lru_counter_1[138] <= 0;lru_counter_2[138] <= 0;tag_1[138] <= 0;tag_2[138] <= 0;cache_mem_1[138] <= 0;cache_mem_2[138] <= 0;
    valid_1[139]  <=   0;valid_2[139]  <=   0;dirty_bit_1[139] <= 0;dirty_bit_2[139] <= 0;lru_counter_1[139] <= 0;lru_counter_2[139] <= 0;tag_1[139] <= 0;tag_2[139] <= 0;cache_mem_1[139] <= 0;cache_mem_2[139] <= 0;
    valid_1[140]  <=   0;valid_2[140]  <=   0;dirty_bit_1[140] <= 0;dirty_bit_2[140] <= 0;lru_counter_1[140] <= 0;lru_counter_2[140] <= 0;tag_1[140] <= 0;tag_2[140] <= 0;cache_mem_1[140] <= 0;cache_mem_2[140] <= 0;
    valid_1[141]  <=   0;valid_2[141]  <=   0;dirty_bit_1[141] <= 0;dirty_bit_2[141] <= 0;lru_counter_1[141] <= 0;lru_counter_2[141] <= 0;tag_1[141] <= 0;tag_2[141] <= 0;cache_mem_1[141] <= 0;cache_mem_2[141] <= 0;
    valid_1[142]  <=   0;valid_2[142]  <=   0;dirty_bit_1[142] <= 0;dirty_bit_2[142] <= 0;lru_counter_1[142] <= 0;lru_counter_2[142] <= 0;tag_1[142] <= 0;tag_2[142] <= 0;cache_mem_1[142] <= 0;cache_mem_2[142] <= 0;
    valid_1[143]  <=   0;valid_2[143]  <=   0;dirty_bit_1[143] <= 0;dirty_bit_2[143] <= 0;lru_counter_1[143] <= 0;lru_counter_2[143] <= 0;tag_1[143] <= 0;tag_2[143] <= 0;cache_mem_1[143] <= 0;cache_mem_2[143] <= 0;
    valid_1[144]  <=   0;valid_2[144]  <=   0;dirty_bit_1[144] <= 0;dirty_bit_2[144] <= 0;lru_counter_1[144] <= 0;lru_counter_2[144] <= 0;tag_1[144] <= 0;tag_2[144] <= 0;cache_mem_1[144] <= 0;cache_mem_2[144] <= 0;
    valid_1[145]  <=   0;valid_2[145]  <=   0;dirty_bit_1[145] <= 0;dirty_bit_2[145] <= 0;lru_counter_1[145] <= 0;lru_counter_2[145] <= 0;tag_1[145] <= 0;tag_2[145] <= 0;cache_mem_1[145] <= 0;cache_mem_2[145] <= 0;
    valid_1[146]  <=   0;valid_2[146]  <=   0;dirty_bit_1[146] <= 0;dirty_bit_2[146] <= 0;lru_counter_1[146] <= 0;lru_counter_2[146] <= 0;tag_1[146] <= 0;tag_2[146] <= 0;cache_mem_1[146] <= 0;cache_mem_2[146] <= 0;
    valid_1[147]  <=   0;valid_2[147]  <=   0;dirty_bit_1[147] <= 0;dirty_bit_2[147] <= 0;lru_counter_1[147] <= 0;lru_counter_2[147] <= 0;tag_1[147] <= 0;tag_2[147] <= 0;cache_mem_1[147] <= 0;cache_mem_2[147] <= 0;
    valid_1[148]  <=   0;valid_2[148]  <=   0;dirty_bit_1[148] <= 0;dirty_bit_2[148] <= 0;lru_counter_1[148] <= 0;lru_counter_2[148] <= 0;tag_1[148] <= 0;tag_2[148] <= 0;cache_mem_1[148] <= 0;cache_mem_2[148] <= 0;
    valid_1[149]  <=   0;valid_2[149]  <=   0;dirty_bit_1[149] <= 0;dirty_bit_2[149] <= 0;lru_counter_1[149] <= 0;lru_counter_2[149] <= 0;tag_1[149] <= 0;tag_2[149] <= 0;cache_mem_1[149] <= 0;cache_mem_2[149] <= 0;
    valid_1[150]  <=   0;valid_2[150]  <=   0;dirty_bit_1[150] <= 0;dirty_bit_2[150] <= 0;lru_counter_1[150] <= 0;lru_counter_2[150] <= 0;tag_1[150] <= 0;tag_2[150] <= 0;cache_mem_1[150] <= 0;cache_mem_2[150] <= 0;
    valid_1[151]  <=   0;valid_2[151]  <=   0;dirty_bit_1[151] <= 0;dirty_bit_2[151] <= 0;lru_counter_1[151] <= 0;lru_counter_2[151] <= 0;tag_1[151] <= 0;tag_2[151] <= 0;cache_mem_1[151] <= 0;cache_mem_2[151] <= 0;
    valid_1[152]  <=   0;valid_2[152]  <=   0;dirty_bit_1[152] <= 0;dirty_bit_2[152] <= 0;lru_counter_1[152] <= 0;lru_counter_2[152] <= 0;tag_1[152] <= 0;tag_2[152] <= 0;cache_mem_1[152] <= 0;cache_mem_2[152] <= 0;
    valid_1[153]  <=   0;valid_2[153]  <=   0;dirty_bit_1[153] <= 0;dirty_bit_2[153] <= 0;lru_counter_1[153] <= 0;lru_counter_2[153] <= 0;tag_1[153] <= 0;tag_2[153] <= 0;cache_mem_1[153] <= 0;cache_mem_2[153] <= 0;
    valid_1[154]  <=   0;valid_2[154]  <=   0;dirty_bit_1[154] <= 0;dirty_bit_2[154] <= 0;lru_counter_1[154] <= 0;lru_counter_2[154] <= 0;tag_1[154] <= 0;tag_2[154] <= 0;cache_mem_1[154] <= 0;cache_mem_2[154] <= 0;
    valid_1[155]  <=   0;valid_2[155]  <=   0;dirty_bit_1[155] <= 0;dirty_bit_2[155] <= 0;lru_counter_1[155] <= 0;lru_counter_2[155] <= 0;tag_1[155] <= 0;tag_2[155] <= 0;cache_mem_1[155] <= 0;cache_mem_2[155] <= 0;
    valid_1[156]  <=   0;valid_2[156]  <=   0;dirty_bit_1[156] <= 0;dirty_bit_2[156] <= 0;lru_counter_1[156] <= 0;lru_counter_2[156] <= 0;tag_1[156] <= 0;tag_2[156] <= 0;cache_mem_1[156] <= 0;cache_mem_2[156] <= 0;
    valid_1[157]  <=   0;valid_2[157]  <=   0;dirty_bit_1[157] <= 0;dirty_bit_2[157] <= 0;lru_counter_1[157] <= 0;lru_counter_2[157] <= 0;tag_1[157] <= 0;tag_2[157] <= 0;cache_mem_1[157] <= 0;cache_mem_2[157] <= 0;
    valid_1[158]  <=   0;valid_2[158]  <=   0;dirty_bit_1[158] <= 0;dirty_bit_2[158] <= 0;lru_counter_1[158] <= 0;lru_counter_2[158] <= 0;tag_1[158] <= 0;tag_2[158] <= 0;cache_mem_1[158] <= 0;cache_mem_2[158] <= 0;
    valid_1[159]  <=   0;valid_2[159]  <=   0;dirty_bit_1[159] <= 0;dirty_bit_2[159] <= 0;lru_counter_1[159] <= 0;lru_counter_2[159] <= 0;tag_1[159] <= 0;tag_2[159] <= 0;cache_mem_1[159] <= 0;cache_mem_2[159] <= 0;
    valid_1[160]  <=   0;valid_2[160]  <=   0;dirty_bit_1[160] <= 0;dirty_bit_2[160] <= 0;lru_counter_1[160] <= 0;lru_counter_2[160] <= 0;tag_1[160] <= 0;tag_2[160] <= 0;cache_mem_1[160] <= 0;cache_mem_2[160] <= 0;
    valid_1[161]  <=   0;valid_2[161]  <=   0;dirty_bit_1[161] <= 0;dirty_bit_2[161] <= 0;lru_counter_1[161] <= 0;lru_counter_2[161] <= 0;tag_1[161] <= 0;tag_2[161] <= 0;cache_mem_1[161] <= 0;cache_mem_2[161] <= 0;
    valid_1[162]  <=   0;valid_2[162]  <=   0;dirty_bit_1[162] <= 0;dirty_bit_2[162] <= 0;lru_counter_1[162] <= 0;lru_counter_2[162] <= 0;tag_1[162] <= 0;tag_2[162] <= 0;cache_mem_1[162] <= 0;cache_mem_2[162] <= 0;
    valid_1[163]  <=   0;valid_2[163]  <=   0;dirty_bit_1[163] <= 0;dirty_bit_2[163] <= 0;lru_counter_1[163] <= 0;lru_counter_2[163] <= 0;tag_1[163] <= 0;tag_2[163] <= 0;cache_mem_1[163] <= 0;cache_mem_2[163] <= 0;
    valid_1[164]  <=   0;valid_2[164]  <=   0;dirty_bit_1[164] <= 0;dirty_bit_2[164] <= 0;lru_counter_1[164] <= 0;lru_counter_2[164] <= 0;tag_1[164] <= 0;tag_2[164] <= 0;cache_mem_1[164] <= 0;cache_mem_2[164] <= 0;
    valid_1[165]  <=   0;valid_2[165]  <=   0;dirty_bit_1[165] <= 0;dirty_bit_2[165] <= 0;lru_counter_1[165] <= 0;lru_counter_2[165] <= 0;tag_1[165] <= 0;tag_2[165] <= 0;cache_mem_1[165] <= 0;cache_mem_2[165] <= 0;
    valid_1[166]  <=   0;valid_2[166]  <=   0;dirty_bit_1[166] <= 0;dirty_bit_2[166] <= 0;lru_counter_1[166] <= 0;lru_counter_2[166] <= 0;tag_1[166] <= 0;tag_2[166] <= 0;cache_mem_1[166] <= 0;cache_mem_2[166] <= 0;
    valid_1[167]  <=   0;valid_2[167]  <=   0;dirty_bit_1[167] <= 0;dirty_bit_2[167] <= 0;lru_counter_1[167] <= 0;lru_counter_2[167] <= 0;tag_1[167] <= 0;tag_2[167] <= 0;cache_mem_1[167] <= 0;cache_mem_2[167] <= 0;
    valid_1[168]  <=   0;valid_2[168]  <=   0;dirty_bit_1[168] <= 0;dirty_bit_2[168] <= 0;lru_counter_1[168] <= 0;lru_counter_2[168] <= 0;tag_1[168] <= 0;tag_2[168] <= 0;cache_mem_1[168] <= 0;cache_mem_2[168] <= 0;
    valid_1[169]  <=   0;valid_2[169]  <=   0;dirty_bit_1[169] <= 0;dirty_bit_2[169] <= 0;lru_counter_1[169] <= 0;lru_counter_2[169] <= 0;tag_1[169] <= 0;tag_2[169] <= 0;cache_mem_1[169] <= 0;cache_mem_2[169] <= 0;
    valid_1[170]  <=   0;valid_2[170]  <=   0;dirty_bit_1[170] <= 0;dirty_bit_2[170] <= 0;lru_counter_1[170] <= 0;lru_counter_2[170] <= 0;tag_1[170] <= 0;tag_2[170] <= 0;cache_mem_1[170] <= 0;cache_mem_2[170] <= 0;
    valid_1[171]  <=   0;valid_2[171]  <=   0;dirty_bit_1[171] <= 0;dirty_bit_2[171] <= 0;lru_counter_1[171] <= 0;lru_counter_2[171] <= 0;tag_1[171] <= 0;tag_2[171] <= 0;cache_mem_1[171] <= 0;cache_mem_2[171] <= 0;
    valid_1[172]  <=   0;valid_2[172]  <=   0;dirty_bit_1[172] <= 0;dirty_bit_2[172] <= 0;lru_counter_1[172] <= 0;lru_counter_2[172] <= 0;tag_1[172] <= 0;tag_2[172] <= 0;cache_mem_1[172] <= 0;cache_mem_2[172] <= 0;
    valid_1[173]  <=   0;valid_2[173]  <=   0;dirty_bit_1[173] <= 0;dirty_bit_2[173] <= 0;lru_counter_1[173] <= 0;lru_counter_2[173] <= 0;tag_1[173] <= 0;tag_2[173] <= 0;cache_mem_1[173] <= 0;cache_mem_2[173] <= 0;
    valid_1[174]  <=   0;valid_2[174]  <=   0;dirty_bit_1[174] <= 0;dirty_bit_2[174] <= 0;lru_counter_1[174] <= 0;lru_counter_2[174] <= 0;tag_1[174] <= 0;tag_2[174] <= 0;cache_mem_1[174] <= 0;cache_mem_2[174] <= 0;
    valid_1[175]  <=   0;valid_2[175]  <=   0;dirty_bit_1[175] <= 0;dirty_bit_2[175] <= 0;lru_counter_1[175] <= 0;lru_counter_2[175] <= 0;tag_1[175] <= 0;tag_2[175] <= 0;cache_mem_1[175] <= 0;cache_mem_2[175] <= 0;
    valid_1[176]  <=   0;valid_2[176]  <=   0;dirty_bit_1[176] <= 0;dirty_bit_2[176] <= 0;lru_counter_1[176] <= 0;lru_counter_2[176] <= 0;tag_1[176] <= 0;tag_2[176] <= 0;cache_mem_1[176] <= 0;cache_mem_2[176] <= 0;
    valid_1[177]  <=   0;valid_2[177]  <=   0;dirty_bit_1[177] <= 0;dirty_bit_2[177] <= 0;lru_counter_1[177] <= 0;lru_counter_2[177] <= 0;tag_1[177] <= 0;tag_2[177] <= 0;cache_mem_1[177] <= 0;cache_mem_2[177] <= 0;
    valid_1[178]  <=   0;valid_2[178]  <=   0;dirty_bit_1[178] <= 0;dirty_bit_2[178] <= 0;lru_counter_1[178] <= 0;lru_counter_2[178] <= 0;tag_1[178] <= 0;tag_2[178] <= 0;cache_mem_1[178] <= 0;cache_mem_2[178] <= 0;
    valid_1[179]  <=   0;valid_2[179]  <=   0;dirty_bit_1[179] <= 0;dirty_bit_2[179] <= 0;lru_counter_1[179] <= 0;lru_counter_2[179] <= 0;tag_1[179] <= 0;tag_2[179] <= 0;cache_mem_1[179] <= 0;cache_mem_2[179] <= 0;
    valid_1[180]  <=   0;valid_2[180]  <=   0;dirty_bit_1[180] <= 0;dirty_bit_2[180] <= 0;lru_counter_1[180] <= 0;lru_counter_2[180] <= 0;tag_1[180] <= 0;tag_2[180] <= 0;cache_mem_1[180] <= 0;cache_mem_2[180] <= 0;
    valid_1[181]  <=   0;valid_2[181]  <=   0;dirty_bit_1[181] <= 0;dirty_bit_2[181] <= 0;lru_counter_1[181] <= 0;lru_counter_2[181] <= 0;tag_1[181] <= 0;tag_2[181] <= 0;cache_mem_1[181] <= 0;cache_mem_2[181] <= 0;
    valid_1[182]  <=   0;valid_2[182]  <=   0;dirty_bit_1[182] <= 0;dirty_bit_2[182] <= 0;lru_counter_1[182] <= 0;lru_counter_2[182] <= 0;tag_1[182] <= 0;tag_2[182] <= 0;cache_mem_1[182] <= 0;cache_mem_2[182] <= 0;
    valid_1[183]  <=   0;valid_2[183]  <=   0;dirty_bit_1[183] <= 0;dirty_bit_2[183] <= 0;lru_counter_1[183] <= 0;lru_counter_2[183] <= 0;tag_1[183] <= 0;tag_2[183] <= 0;cache_mem_1[183] <= 0;cache_mem_2[183] <= 0;
    valid_1[184]  <=   0;valid_2[184]  <=   0;dirty_bit_1[184] <= 0;dirty_bit_2[184] <= 0;lru_counter_1[184] <= 0;lru_counter_2[184] <= 0;tag_1[184] <= 0;tag_2[184] <= 0;cache_mem_1[184] <= 0;cache_mem_2[184] <= 0;
    valid_1[185]  <=   0;valid_2[185]  <=   0;dirty_bit_1[185] <= 0;dirty_bit_2[185] <= 0;lru_counter_1[185] <= 0;lru_counter_2[185] <= 0;tag_1[185] <= 0;tag_2[185] <= 0;cache_mem_1[185] <= 0;cache_mem_2[185] <= 0;
    valid_1[186]  <=   0;valid_2[186]  <=   0;dirty_bit_1[186] <= 0;dirty_bit_2[186] <= 0;lru_counter_1[186] <= 0;lru_counter_2[186] <= 0;tag_1[186] <= 0;tag_2[186] <= 0;cache_mem_1[186] <= 0;cache_mem_2[186] <= 0;
    valid_1[187]  <=   0;valid_2[187]  <=   0;dirty_bit_1[187] <= 0;dirty_bit_2[187] <= 0;lru_counter_1[187] <= 0;lru_counter_2[187] <= 0;tag_1[187] <= 0;tag_2[187] <= 0;cache_mem_1[187] <= 0;cache_mem_2[187] <= 0;
    valid_1[188]  <=   0;valid_2[188]  <=   0;dirty_bit_1[188] <= 0;dirty_bit_2[188] <= 0;lru_counter_1[188] <= 0;lru_counter_2[188] <= 0;tag_1[188] <= 0;tag_2[188] <= 0;cache_mem_1[188] <= 0;cache_mem_2[188] <= 0;
    valid_1[189]  <=   0;valid_2[189]  <=   0;dirty_bit_1[189] <= 0;dirty_bit_2[189] <= 0;lru_counter_1[189] <= 0;lru_counter_2[189] <= 0;tag_1[189] <= 0;tag_2[189] <= 0;cache_mem_1[189] <= 0;cache_mem_2[189] <= 0;
    valid_1[190]  <=   0;valid_2[190]  <=   0;dirty_bit_1[190] <= 0;dirty_bit_2[190] <= 0;lru_counter_1[190] <= 0;lru_counter_2[190] <= 0;tag_1[190] <= 0;tag_2[190] <= 0;cache_mem_1[190] <= 0;cache_mem_2[190] <= 0;
    valid_1[191]  <=   0;valid_2[191]  <=   0;dirty_bit_1[191] <= 0;dirty_bit_2[191] <= 0;lru_counter_1[191] <= 0;lru_counter_2[191] <= 0;tag_1[191] <= 0;tag_2[191] <= 0;cache_mem_1[191] <= 0;cache_mem_2[191] <= 0;
    valid_1[192]  <=   0;valid_2[192]  <=   0;dirty_bit_1[192] <= 0;dirty_bit_2[192] <= 0;lru_counter_1[192] <= 0;lru_counter_2[192] <= 0;tag_1[192] <= 0;tag_2[192] <= 0;cache_mem_1[192] <= 0;cache_mem_2[192] <= 0;
    valid_1[193]  <=   0;valid_2[193]  <=   0;dirty_bit_1[193] <= 0;dirty_bit_2[193] <= 0;lru_counter_1[193] <= 0;lru_counter_2[193] <= 0;tag_1[193] <= 0;tag_2[193] <= 0;cache_mem_1[193] <= 0;cache_mem_2[193] <= 0;
    valid_1[194]  <=   0;valid_2[194]  <=   0;dirty_bit_1[194] <= 0;dirty_bit_2[194] <= 0;lru_counter_1[194] <= 0;lru_counter_2[194] <= 0;tag_1[194] <= 0;tag_2[194] <= 0;cache_mem_1[194] <= 0;cache_mem_2[194] <= 0;
    valid_1[195]  <=   0;valid_2[195]  <=   0;dirty_bit_1[195] <= 0;dirty_bit_2[195] <= 0;lru_counter_1[195] <= 0;lru_counter_2[195] <= 0;tag_1[195] <= 0;tag_2[195] <= 0;cache_mem_1[195] <= 0;cache_mem_2[195] <= 0;
    valid_1[196]  <=   0;valid_2[196]  <=   0;dirty_bit_1[196] <= 0;dirty_bit_2[196] <= 0;lru_counter_1[196] <= 0;lru_counter_2[196] <= 0;tag_1[196] <= 0;tag_2[196] <= 0;cache_mem_1[196] <= 0;cache_mem_2[196] <= 0;
    valid_1[197]  <=   0;valid_2[197]  <=   0;dirty_bit_1[197] <= 0;dirty_bit_2[197] <= 0;lru_counter_1[197] <= 0;lru_counter_2[197] <= 0;tag_1[197] <= 0;tag_2[197] <= 0;cache_mem_1[197] <= 0;cache_mem_2[197] <= 0;
    valid_1[198]  <=   0;valid_2[198]  <=   0;dirty_bit_1[198] <= 0;dirty_bit_2[198] <= 0;lru_counter_1[198] <= 0;lru_counter_2[198] <= 0;tag_1[198] <= 0;tag_2[198] <= 0;cache_mem_1[198] <= 0;cache_mem_2[198] <= 0;
    valid_1[199]  <=   0;valid_2[199]  <=   0;dirty_bit_1[199] <= 0;dirty_bit_2[199] <= 0;lru_counter_1[199] <= 0;lru_counter_2[199] <= 0;tag_1[199] <= 0;tag_2[199] <= 0;cache_mem_1[199] <= 0;cache_mem_2[199] <= 0;
    valid_1[200]  <=   0;valid_2[200]  <=   0;dirty_bit_1[200] <= 0;dirty_bit_2[200] <= 0;lru_counter_1[200] <= 0;lru_counter_2[200] <= 0;tag_1[200] <= 0;tag_2[200] <= 0;cache_mem_1[200] <= 0;cache_mem_2[200] <= 0;
    valid_1[201]  <=   0;valid_2[201]  <=   0;dirty_bit_1[201] <= 0;dirty_bit_2[201] <= 0;lru_counter_1[201] <= 0;lru_counter_2[201] <= 0;tag_1[201] <= 0;tag_2[201] <= 0;cache_mem_1[201] <= 0;cache_mem_2[201] <= 0;
    valid_1[202]  <=   0;valid_2[202]  <=   0;dirty_bit_1[202] <= 0;dirty_bit_2[202] <= 0;lru_counter_1[202] <= 0;lru_counter_2[202] <= 0;tag_1[202] <= 0;tag_2[202] <= 0;cache_mem_1[202] <= 0;cache_mem_2[202] <= 0;
    valid_1[203]  <=   0;valid_2[203]  <=   0;dirty_bit_1[203] <= 0;dirty_bit_2[203] <= 0;lru_counter_1[203] <= 0;lru_counter_2[203] <= 0;tag_1[203] <= 0;tag_2[203] <= 0;cache_mem_1[203] <= 0;cache_mem_2[203] <= 0;
    valid_1[204]  <=   0;valid_2[204]  <=   0;dirty_bit_1[204] <= 0;dirty_bit_2[204] <= 0;lru_counter_1[204] <= 0;lru_counter_2[204] <= 0;tag_1[204] <= 0;tag_2[204] <= 0;cache_mem_1[204] <= 0;cache_mem_2[204] <= 0;
    valid_1[205]  <=   0;valid_2[205]  <=   0;dirty_bit_1[205] <= 0;dirty_bit_2[205] <= 0;lru_counter_1[205] <= 0;lru_counter_2[205] <= 0;tag_1[205] <= 0;tag_2[205] <= 0;cache_mem_1[205] <= 0;cache_mem_2[205] <= 0;
    valid_1[206]  <=   0;valid_2[206]  <=   0;dirty_bit_1[206] <= 0;dirty_bit_2[206] <= 0;lru_counter_1[206] <= 0;lru_counter_2[206] <= 0;tag_1[206] <= 0;tag_2[206] <= 0;cache_mem_1[206] <= 0;cache_mem_2[206] <= 0;
    valid_1[207]  <=   0;valid_2[207]  <=   0;dirty_bit_1[207] <= 0;dirty_bit_2[207] <= 0;lru_counter_1[207] <= 0;lru_counter_2[207] <= 0;tag_1[207] <= 0;tag_2[207] <= 0;cache_mem_1[207] <= 0;cache_mem_2[207] <= 0;
    valid_1[208]  <=   0;valid_2[208]  <=   0;dirty_bit_1[208] <= 0;dirty_bit_2[208] <= 0;lru_counter_1[208] <= 0;lru_counter_2[208] <= 0;tag_1[208] <= 0;tag_2[208] <= 0;cache_mem_1[208] <= 0;cache_mem_2[208] <= 0;
    valid_1[209]  <=   0;valid_2[209]  <=   0;dirty_bit_1[209] <= 0;dirty_bit_2[209] <= 0;lru_counter_1[209] <= 0;lru_counter_2[209] <= 0;tag_1[209] <= 0;tag_2[209] <= 0;cache_mem_1[209] <= 0;cache_mem_2[209] <= 0;
    valid_1[210]  <=   0;valid_2[210]  <=   0;dirty_bit_1[210] <= 0;dirty_bit_2[210] <= 0;lru_counter_1[210] <= 0;lru_counter_2[210] <= 0;tag_1[210] <= 0;tag_2[210] <= 0;cache_mem_1[210] <= 0;cache_mem_2[210] <= 0;
    valid_1[211]  <=   0;valid_2[211]  <=   0;dirty_bit_1[211] <= 0;dirty_bit_2[211] <= 0;lru_counter_1[211] <= 0;lru_counter_2[211] <= 0;tag_1[211] <= 0;tag_2[211] <= 0;cache_mem_1[211] <= 0;cache_mem_2[211] <= 0;
    valid_1[212]  <=   0;valid_2[212]  <=   0;dirty_bit_1[212] <= 0;dirty_bit_2[212] <= 0;lru_counter_1[212] <= 0;lru_counter_2[212] <= 0;tag_1[212] <= 0;tag_2[212] <= 0;cache_mem_1[212] <= 0;cache_mem_2[212] <= 0;
    valid_1[213]  <=   0;valid_2[213]  <=   0;dirty_bit_1[213] <= 0;dirty_bit_2[213] <= 0;lru_counter_1[213] <= 0;lru_counter_2[213] <= 0;tag_1[213] <= 0;tag_2[213] <= 0;cache_mem_1[213] <= 0;cache_mem_2[213] <= 0;
    valid_1[214]  <=   0;valid_2[214]  <=   0;dirty_bit_1[214] <= 0;dirty_bit_2[214] <= 0;lru_counter_1[214] <= 0;lru_counter_2[214] <= 0;tag_1[214] <= 0;tag_2[214] <= 0;cache_mem_1[214] <= 0;cache_mem_2[214] <= 0;
    valid_1[215]  <=   0;valid_2[215]  <=   0;dirty_bit_1[215] <= 0;dirty_bit_2[215] <= 0;lru_counter_1[215] <= 0;lru_counter_2[215] <= 0;tag_1[215] <= 0;tag_2[215] <= 0;cache_mem_1[215] <= 0;cache_mem_2[215] <= 0;
    valid_1[216]  <=   0;valid_2[216]  <=   0;dirty_bit_1[216] <= 0;dirty_bit_2[216] <= 0;lru_counter_1[216] <= 0;lru_counter_2[216] <= 0;tag_1[216] <= 0;tag_2[216] <= 0;cache_mem_1[216] <= 0;cache_mem_2[216] <= 0;
    valid_1[217]  <=   0;valid_2[217]  <=   0;dirty_bit_1[217] <= 0;dirty_bit_2[217] <= 0;lru_counter_1[217] <= 0;lru_counter_2[217] <= 0;tag_1[217] <= 0;tag_2[217] <= 0;cache_mem_1[217] <= 0;cache_mem_2[217] <= 0;
    valid_1[218]  <=   0;valid_2[218]  <=   0;dirty_bit_1[218] <= 0;dirty_bit_2[218] <= 0;lru_counter_1[218] <= 0;lru_counter_2[218] <= 0;tag_1[218] <= 0;tag_2[218] <= 0;cache_mem_1[218] <= 0;cache_mem_2[218] <= 0;
    valid_1[219]  <=   0;valid_2[219]  <=   0;dirty_bit_1[219] <= 0;dirty_bit_2[219] <= 0;lru_counter_1[219] <= 0;lru_counter_2[219] <= 0;tag_1[219] <= 0;tag_2[219] <= 0;cache_mem_1[219] <= 0;cache_mem_2[219] <= 0;
    valid_1[220]  <=   0;valid_2[220]  <=   0;dirty_bit_1[220] <= 0;dirty_bit_2[220] <= 0;lru_counter_1[220] <= 0;lru_counter_2[220] <= 0;tag_1[220] <= 0;tag_2[220] <= 0;cache_mem_1[220] <= 0;cache_mem_2[220] <= 0;
    valid_1[221]  <=   0;valid_2[221]  <=   0;dirty_bit_1[221] <= 0;dirty_bit_2[221] <= 0;lru_counter_1[221] <= 0;lru_counter_2[221] <= 0;tag_1[221] <= 0;tag_2[221] <= 0;cache_mem_1[221] <= 0;cache_mem_2[221] <= 0;
    valid_1[222]  <=   0;valid_2[222]  <=   0;dirty_bit_1[222] <= 0;dirty_bit_2[222] <= 0;lru_counter_1[222] <= 0;lru_counter_2[222] <= 0;tag_1[222] <= 0;tag_2[222] <= 0;cache_mem_1[222] <= 0;cache_mem_2[222] <= 0;
    valid_1[223]  <=   0;valid_2[223]  <=   0;dirty_bit_1[223] <= 0;dirty_bit_2[223] <= 0;lru_counter_1[223] <= 0;lru_counter_2[223] <= 0;tag_1[223] <= 0;tag_2[223] <= 0;cache_mem_1[223] <= 0;cache_mem_2[223] <= 0;
    valid_1[224]  <=   0;valid_2[224]  <=   0;dirty_bit_1[224] <= 0;dirty_bit_2[224] <= 0;lru_counter_1[224] <= 0;lru_counter_2[224] <= 0;tag_1[224] <= 0;tag_2[224] <= 0;cache_mem_1[224] <= 0;cache_mem_2[224] <= 0;
    valid_1[225]  <=   0;valid_2[225]  <=   0;dirty_bit_1[225] <= 0;dirty_bit_2[225] <= 0;lru_counter_1[225] <= 0;lru_counter_2[225] <= 0;tag_1[225] <= 0;tag_2[225] <= 0;cache_mem_1[225] <= 0;cache_mem_2[225] <= 0;
    valid_1[226]  <=   0;valid_2[226]  <=   0;dirty_bit_1[226] <= 0;dirty_bit_2[226] <= 0;lru_counter_1[226] <= 0;lru_counter_2[226] <= 0;tag_1[226] <= 0;tag_2[226] <= 0;cache_mem_1[226] <= 0;cache_mem_2[226] <= 0;
    valid_1[227]  <=   0;valid_2[227]  <=   0;dirty_bit_1[227] <= 0;dirty_bit_2[227] <= 0;lru_counter_1[227] <= 0;lru_counter_2[227] <= 0;tag_1[227] <= 0;tag_2[227] <= 0;cache_mem_1[227] <= 0;cache_mem_2[227] <= 0;
    valid_1[228]  <=   0;valid_2[228]  <=   0;dirty_bit_1[228] <= 0;dirty_bit_2[228] <= 0;lru_counter_1[228] <= 0;lru_counter_2[228] <= 0;tag_1[228] <= 0;tag_2[228] <= 0;cache_mem_1[228] <= 0;cache_mem_2[228] <= 0;
    valid_1[229]  <=   0;valid_2[229]  <=   0;dirty_bit_1[229] <= 0;dirty_bit_2[229] <= 0;lru_counter_1[229] <= 0;lru_counter_2[229] <= 0;tag_1[229] <= 0;tag_2[229] <= 0;cache_mem_1[229] <= 0;cache_mem_2[229] <= 0;
    valid_1[230]  <=   0;valid_2[230]  <=   0;dirty_bit_1[230] <= 0;dirty_bit_2[230] <= 0;lru_counter_1[230] <= 0;lru_counter_2[230] <= 0;tag_1[230] <= 0;tag_2[230] <= 0;cache_mem_1[230] <= 0;cache_mem_2[230] <= 0;
    valid_1[231]  <=   0;valid_2[231]  <=   0;dirty_bit_1[231] <= 0;dirty_bit_2[231] <= 0;lru_counter_1[231] <= 0;lru_counter_2[231] <= 0;tag_1[231] <= 0;tag_2[231] <= 0;cache_mem_1[231] <= 0;cache_mem_2[231] <= 0;
    valid_1[232]  <=   0;valid_2[232]  <=   0;dirty_bit_1[232] <= 0;dirty_bit_2[232] <= 0;lru_counter_1[232] <= 0;lru_counter_2[232] <= 0;tag_1[232] <= 0;tag_2[232] <= 0;cache_mem_1[232] <= 0;cache_mem_2[232] <= 0;
    valid_1[233]  <=   0;valid_2[233]  <=   0;dirty_bit_1[233] <= 0;dirty_bit_2[233] <= 0;lru_counter_1[233] <= 0;lru_counter_2[233] <= 0;tag_1[233] <= 0;tag_2[233] <= 0;cache_mem_1[233] <= 0;cache_mem_2[233] <= 0;
    valid_1[234]  <=   0;valid_2[234]  <=   0;dirty_bit_1[234] <= 0;dirty_bit_2[234] <= 0;lru_counter_1[234] <= 0;lru_counter_2[234] <= 0;tag_1[234] <= 0;tag_2[234] <= 0;cache_mem_1[234] <= 0;cache_mem_2[234] <= 0;
    valid_1[235]  <=   0;valid_2[235]  <=   0;dirty_bit_1[235] <= 0;dirty_bit_2[235] <= 0;lru_counter_1[235] <= 0;lru_counter_2[235] <= 0;tag_1[235] <= 0;tag_2[235] <= 0;cache_mem_1[235] <= 0;cache_mem_2[235] <= 0;
    valid_1[236]  <=   0;valid_2[236]  <=   0;dirty_bit_1[236] <= 0;dirty_bit_2[236] <= 0;lru_counter_1[236] <= 0;lru_counter_2[236] <= 0;tag_1[236] <= 0;tag_2[236] <= 0;cache_mem_1[236] <= 0;cache_mem_2[236] <= 0;
    valid_1[237]  <=   0;valid_2[237]  <=   0;dirty_bit_1[237] <= 0;dirty_bit_2[237] <= 0;lru_counter_1[237] <= 0;lru_counter_2[237] <= 0;tag_1[237] <= 0;tag_2[237] <= 0;cache_mem_1[237] <= 0;cache_mem_2[237] <= 0;
    valid_1[238]  <=   0;valid_2[238]  <=   0;dirty_bit_1[238] <= 0;dirty_bit_2[238] <= 0;lru_counter_1[238] <= 0;lru_counter_2[238] <= 0;tag_1[238] <= 0;tag_2[238] <= 0;cache_mem_1[238] <= 0;cache_mem_2[238] <= 0;
    valid_1[239]  <=   0;valid_2[239]  <=   0;dirty_bit_1[239] <= 0;dirty_bit_2[239] <= 0;lru_counter_1[239] <= 0;lru_counter_2[239] <= 0;tag_1[239] <= 0;tag_2[239] <= 0;cache_mem_1[239] <= 0;cache_mem_2[239] <= 0;
    valid_1[240]  <=   0;valid_2[240]  <=   0;dirty_bit_1[240] <= 0;dirty_bit_2[240] <= 0;lru_counter_1[240] <= 0;lru_counter_2[240] <= 0;tag_1[240] <= 0;tag_2[240] <= 0;cache_mem_1[240] <= 0;cache_mem_2[240] <= 0;
    valid_1[241]  <=   0;valid_2[241]  <=   0;dirty_bit_1[241] <= 0;dirty_bit_2[241] <= 0;lru_counter_1[241] <= 0;lru_counter_2[241] <= 0;tag_1[241] <= 0;tag_2[241] <= 0;cache_mem_1[241] <= 0;cache_mem_2[241] <= 0;
    valid_1[242]  <=   0;valid_2[242]  <=   0;dirty_bit_1[242] <= 0;dirty_bit_2[242] <= 0;lru_counter_1[242] <= 0;lru_counter_2[242] <= 0;tag_1[242] <= 0;tag_2[242] <= 0;cache_mem_1[242] <= 0;cache_mem_2[242] <= 0;
    valid_1[243]  <=   0;valid_2[243]  <=   0;dirty_bit_1[243] <= 0;dirty_bit_2[243] <= 0;lru_counter_1[243] <= 0;lru_counter_2[243] <= 0;tag_1[243] <= 0;tag_2[243] <= 0;cache_mem_1[243] <= 0;cache_mem_2[243] <= 0;
    valid_1[244]  <=   0;valid_2[244]  <=   0;dirty_bit_1[244] <= 0;dirty_bit_2[244] <= 0;lru_counter_1[244] <= 0;lru_counter_2[244] <= 0;tag_1[244] <= 0;tag_2[244] <= 0;cache_mem_1[244] <= 0;cache_mem_2[244] <= 0;
    valid_1[245]  <=   0;valid_2[245]  <=   0;dirty_bit_1[245] <= 0;dirty_bit_2[245] <= 0;lru_counter_1[245] <= 0;lru_counter_2[245] <= 0;tag_1[245] <= 0;tag_2[245] <= 0;cache_mem_1[245] <= 0;cache_mem_2[245] <= 0;
    valid_1[246]  <=   0;valid_2[246]  <=   0;dirty_bit_1[246] <= 0;dirty_bit_2[246] <= 0;lru_counter_1[246] <= 0;lru_counter_2[246] <= 0;tag_1[246] <= 0;tag_2[246] <= 0;cache_mem_1[246] <= 0;cache_mem_2[246] <= 0;
    valid_1[247]  <=   0;valid_2[247]  <=   0;dirty_bit_1[247] <= 0;dirty_bit_2[247] <= 0;lru_counter_1[247] <= 0;lru_counter_2[247] <= 0;tag_1[247] <= 0;tag_2[247] <= 0;cache_mem_1[247] <= 0;cache_mem_2[247] <= 0;
    valid_1[248]  <=   0;valid_2[248]  <=   0;dirty_bit_1[248] <= 0;dirty_bit_2[248] <= 0;lru_counter_1[248] <= 0;lru_counter_2[248] <= 0;tag_1[248] <= 0;tag_2[248] <= 0;cache_mem_1[248] <= 0;cache_mem_2[248] <= 0;
    valid_1[249]  <=   0;valid_2[249]  <=   0;dirty_bit_1[249] <= 0;dirty_bit_2[249] <= 0;lru_counter_1[249] <= 0;lru_counter_2[249] <= 0;tag_1[249] <= 0;tag_2[249] <= 0;cache_mem_1[249] <= 0;cache_mem_2[249] <= 0;
    valid_1[250]  <=   0;valid_2[250]  <=   0;dirty_bit_1[250] <= 0;dirty_bit_2[250] <= 0;lru_counter_1[250] <= 0;lru_counter_2[250] <= 0;tag_1[250] <= 0;tag_2[250] <= 0;cache_mem_1[250] <= 0;cache_mem_2[250] <= 0;
    valid_1[251]  <=   0;valid_2[251]  <=   0;dirty_bit_1[251] <= 0;dirty_bit_2[251] <= 0;lru_counter_1[251] <= 0;lru_counter_2[251] <= 0;tag_1[251] <= 0;tag_2[251] <= 0;cache_mem_1[251] <= 0;cache_mem_2[251] <= 0;
    valid_1[252]  <=   0;valid_2[252]  <=   0;dirty_bit_1[252] <= 0;dirty_bit_2[252] <= 0;lru_counter_1[252] <= 0;lru_counter_2[252] <= 0;tag_1[252] <= 0;tag_2[252] <= 0;cache_mem_1[252] <= 0;cache_mem_2[252] <= 0;
    valid_1[253]  <=   0;valid_2[253]  <=   0;dirty_bit_1[253] <= 0;dirty_bit_2[253] <= 0;lru_counter_1[253] <= 0;lru_counter_2[253] <= 0;tag_1[253] <= 0;tag_2[253] <= 0;cache_mem_1[253] <= 0;cache_mem_2[253] <= 0;
    valid_1[254]  <=   0;valid_2[254]  <=   0;dirty_bit_1[254] <= 0;dirty_bit_2[254] <= 0;lru_counter_1[254] <= 0;lru_counter_2[254] <= 0;tag_1[254] <= 0;tag_2[254] <= 0;cache_mem_1[254] <= 0;cache_mem_2[254] <= 0;
    valid_1[255]  <=   0;valid_2[255]  <=   0;dirty_bit_1[255] <= 0;dirty_bit_2[255] <= 0;lru_counter_1[255] <= 0;lru_counter_2[255] <= 0;tag_1[255] <= 0;tag_2[255] <= 0;cache_mem_1[255] <= 0;cache_mem_2[255] <= 0;
    valid_1[256]  <=   0;valid_2[256]  <=   0;dirty_bit_1[256] <= 0;dirty_bit_2[256] <= 0;lru_counter_1[256] <= 0;lru_counter_2[256] <= 0;tag_1[256] <= 0;tag_2[256] <= 0;cache_mem_1[256] <= 0;cache_mem_2[256] <= 0;
    valid_1[257]  <=   0;valid_2[257]  <=   0;dirty_bit_1[257] <= 0;dirty_bit_2[257] <= 0;lru_counter_1[257] <= 0;lru_counter_2[257] <= 0;tag_1[257] <= 0;tag_2[257] <= 0;cache_mem_1[257] <= 0;cache_mem_2[257] <= 0;
    valid_1[258]  <=   0;valid_2[258]  <=   0;dirty_bit_1[258] <= 0;dirty_bit_2[258] <= 0;lru_counter_1[258] <= 0;lru_counter_2[258] <= 0;tag_1[258] <= 0;tag_2[258] <= 0;cache_mem_1[258] <= 0;cache_mem_2[258] <= 0;
    valid_1[259]  <=   0;valid_2[259]  <=   0;dirty_bit_1[259] <= 0;dirty_bit_2[259] <= 0;lru_counter_1[259] <= 0;lru_counter_2[259] <= 0;tag_1[259] <= 0;tag_2[259] <= 0;cache_mem_1[259] <= 0;cache_mem_2[259] <= 0;
    valid_1[260]  <=   0;valid_2[260]  <=   0;dirty_bit_1[260] <= 0;dirty_bit_2[260] <= 0;lru_counter_1[260] <= 0;lru_counter_2[260] <= 0;tag_1[260] <= 0;tag_2[260] <= 0;cache_mem_1[260] <= 0;cache_mem_2[260] <= 0;
    valid_1[261]  <=   0;valid_2[261]  <=   0;dirty_bit_1[261] <= 0;dirty_bit_2[261] <= 0;lru_counter_1[261] <= 0;lru_counter_2[261] <= 0;tag_1[261] <= 0;tag_2[261] <= 0;cache_mem_1[261] <= 0;cache_mem_2[261] <= 0;
    valid_1[262]  <=   0;valid_2[262]  <=   0;dirty_bit_1[262] <= 0;dirty_bit_2[262] <= 0;lru_counter_1[262] <= 0;lru_counter_2[262] <= 0;tag_1[262] <= 0;tag_2[262] <= 0;cache_mem_1[262] <= 0;cache_mem_2[262] <= 0;
    valid_1[263]  <=   0;valid_2[263]  <=   0;dirty_bit_1[263] <= 0;dirty_bit_2[263] <= 0;lru_counter_1[263] <= 0;lru_counter_2[263] <= 0;tag_1[263] <= 0;tag_2[263] <= 0;cache_mem_1[263] <= 0;cache_mem_2[263] <= 0;
    valid_1[264]  <=   0;valid_2[264]  <=   0;dirty_bit_1[264] <= 0;dirty_bit_2[264] <= 0;lru_counter_1[264] <= 0;lru_counter_2[264] <= 0;tag_1[264] <= 0;tag_2[264] <= 0;cache_mem_1[264] <= 0;cache_mem_2[264] <= 0;
    valid_1[265]  <=   0;valid_2[265]  <=   0;dirty_bit_1[265] <= 0;dirty_bit_2[265] <= 0;lru_counter_1[265] <= 0;lru_counter_2[265] <= 0;tag_1[265] <= 0;tag_2[265] <= 0;cache_mem_1[265] <= 0;cache_mem_2[265] <= 0;
    valid_1[266]  <=   0;valid_2[266]  <=   0;dirty_bit_1[266] <= 0;dirty_bit_2[266] <= 0;lru_counter_1[266] <= 0;lru_counter_2[266] <= 0;tag_1[266] <= 0;tag_2[266] <= 0;cache_mem_1[266] <= 0;cache_mem_2[266] <= 0;
    valid_1[267]  <=   0;valid_2[267]  <=   0;dirty_bit_1[267] <= 0;dirty_bit_2[267] <= 0;lru_counter_1[267] <= 0;lru_counter_2[267] <= 0;tag_1[267] <= 0;tag_2[267] <= 0;cache_mem_1[267] <= 0;cache_mem_2[267] <= 0;
    valid_1[268]  <=   0;valid_2[268]  <=   0;dirty_bit_1[268] <= 0;dirty_bit_2[268] <= 0;lru_counter_1[268] <= 0;lru_counter_2[268] <= 0;tag_1[268] <= 0;tag_2[268] <= 0;cache_mem_1[268] <= 0;cache_mem_2[268] <= 0;
    valid_1[269]  <=   0;valid_2[269]  <=   0;dirty_bit_1[269] <= 0;dirty_bit_2[269] <= 0;lru_counter_1[269] <= 0;lru_counter_2[269] <= 0;tag_1[269] <= 0;tag_2[269] <= 0;cache_mem_1[269] <= 0;cache_mem_2[269] <= 0;
    valid_1[270]  <=   0;valid_2[270]  <=   0;dirty_bit_1[270] <= 0;dirty_bit_2[270] <= 0;lru_counter_1[270] <= 0;lru_counter_2[270] <= 0;tag_1[270] <= 0;tag_2[270] <= 0;cache_mem_1[270] <= 0;cache_mem_2[270] <= 0;
    valid_1[271]  <=   0;valid_2[271]  <=   0;dirty_bit_1[271] <= 0;dirty_bit_2[271] <= 0;lru_counter_1[271] <= 0;lru_counter_2[271] <= 0;tag_1[271] <= 0;tag_2[271] <= 0;cache_mem_1[271] <= 0;cache_mem_2[271] <= 0;
    valid_1[272]  <=   0;valid_2[272]  <=   0;dirty_bit_1[272] <= 0;dirty_bit_2[272] <= 0;lru_counter_1[272] <= 0;lru_counter_2[272] <= 0;tag_1[272] <= 0;tag_2[272] <= 0;cache_mem_1[272] <= 0;cache_mem_2[272] <= 0;
    valid_1[273]  <=   0;valid_2[273]  <=   0;dirty_bit_1[273] <= 0;dirty_bit_2[273] <= 0;lru_counter_1[273] <= 0;lru_counter_2[273] <= 0;tag_1[273] <= 0;tag_2[273] <= 0;cache_mem_1[273] <= 0;cache_mem_2[273] <= 0;
    valid_1[274]  <=   0;valid_2[274]  <=   0;dirty_bit_1[274] <= 0;dirty_bit_2[274] <= 0;lru_counter_1[274] <= 0;lru_counter_2[274] <= 0;tag_1[274] <= 0;tag_2[274] <= 0;cache_mem_1[274] <= 0;cache_mem_2[274] <= 0;
    valid_1[275]  <=   0;valid_2[275]  <=   0;dirty_bit_1[275] <= 0;dirty_bit_2[275] <= 0;lru_counter_1[275] <= 0;lru_counter_2[275] <= 0;tag_1[275] <= 0;tag_2[275] <= 0;cache_mem_1[275] <= 0;cache_mem_2[275] <= 0;
    valid_1[276]  <=   0;valid_2[276]  <=   0;dirty_bit_1[276] <= 0;dirty_bit_2[276] <= 0;lru_counter_1[276] <= 0;lru_counter_2[276] <= 0;tag_1[276] <= 0;tag_2[276] <= 0;cache_mem_1[276] <= 0;cache_mem_2[276] <= 0;
    valid_1[277]  <=   0;valid_2[277]  <=   0;dirty_bit_1[277] <= 0;dirty_bit_2[277] <= 0;lru_counter_1[277] <= 0;lru_counter_2[277] <= 0;tag_1[277] <= 0;tag_2[277] <= 0;cache_mem_1[277] <= 0;cache_mem_2[277] <= 0;
    valid_1[278]  <=   0;valid_2[278]  <=   0;dirty_bit_1[278] <= 0;dirty_bit_2[278] <= 0;lru_counter_1[278] <= 0;lru_counter_2[278] <= 0;tag_1[278] <= 0;tag_2[278] <= 0;cache_mem_1[278] <= 0;cache_mem_2[278] <= 0;
    valid_1[279]  <=   0;valid_2[279]  <=   0;dirty_bit_1[279] <= 0;dirty_bit_2[279] <= 0;lru_counter_1[279] <= 0;lru_counter_2[279] <= 0;tag_1[279] <= 0;tag_2[279] <= 0;cache_mem_1[279] <= 0;cache_mem_2[279] <= 0;
    valid_1[280]  <=   0;valid_2[280]  <=   0;dirty_bit_1[280] <= 0;dirty_bit_2[280] <= 0;lru_counter_1[280] <= 0;lru_counter_2[280] <= 0;tag_1[280] <= 0;tag_2[280] <= 0;cache_mem_1[280] <= 0;cache_mem_2[280] <= 0;
    valid_1[281]  <=   0;valid_2[281]  <=   0;dirty_bit_1[281] <= 0;dirty_bit_2[281] <= 0;lru_counter_1[281] <= 0;lru_counter_2[281] <= 0;tag_1[281] <= 0;tag_2[281] <= 0;cache_mem_1[281] <= 0;cache_mem_2[281] <= 0;
    valid_1[282]  <=   0;valid_2[282]  <=   0;dirty_bit_1[282] <= 0;dirty_bit_2[282] <= 0;lru_counter_1[282] <= 0;lru_counter_2[282] <= 0;tag_1[282] <= 0;tag_2[282] <= 0;cache_mem_1[282] <= 0;cache_mem_2[282] <= 0;
    valid_1[283]  <=   0;valid_2[283]  <=   0;dirty_bit_1[283] <= 0;dirty_bit_2[283] <= 0;lru_counter_1[283] <= 0;lru_counter_2[283] <= 0;tag_1[283] <= 0;tag_2[283] <= 0;cache_mem_1[283] <= 0;cache_mem_2[283] <= 0;
    valid_1[284]  <=   0;valid_2[284]  <=   0;dirty_bit_1[284] <= 0;dirty_bit_2[284] <= 0;lru_counter_1[284] <= 0;lru_counter_2[284] <= 0;tag_1[284] <= 0;tag_2[284] <= 0;cache_mem_1[284] <= 0;cache_mem_2[284] <= 0;
    valid_1[285]  <=   0;valid_2[285]  <=   0;dirty_bit_1[285] <= 0;dirty_bit_2[285] <= 0;lru_counter_1[285] <= 0;lru_counter_2[285] <= 0;tag_1[285] <= 0;tag_2[285] <= 0;cache_mem_1[285] <= 0;cache_mem_2[285] <= 0;
    valid_1[286]  <=   0;valid_2[286]  <=   0;dirty_bit_1[286] <= 0;dirty_bit_2[286] <= 0;lru_counter_1[286] <= 0;lru_counter_2[286] <= 0;tag_1[286] <= 0;tag_2[286] <= 0;cache_mem_1[286] <= 0;cache_mem_2[286] <= 0;
    valid_1[287]  <=   0;valid_2[287]  <=   0;dirty_bit_1[287] <= 0;dirty_bit_2[287] <= 0;lru_counter_1[287] <= 0;lru_counter_2[287] <= 0;tag_1[287] <= 0;tag_2[287] <= 0;cache_mem_1[287] <= 0;cache_mem_2[287] <= 0;
    valid_1[288]  <=   0;valid_2[288]  <=   0;dirty_bit_1[288] <= 0;dirty_bit_2[288] <= 0;lru_counter_1[288] <= 0;lru_counter_2[288] <= 0;tag_1[288] <= 0;tag_2[288] <= 0;cache_mem_1[288] <= 0;cache_mem_2[288] <= 0;
    valid_1[289]  <=   0;valid_2[289]  <=   0;dirty_bit_1[289] <= 0;dirty_bit_2[289] <= 0;lru_counter_1[289] <= 0;lru_counter_2[289] <= 0;tag_1[289] <= 0;tag_2[289] <= 0;cache_mem_1[289] <= 0;cache_mem_2[289] <= 0;
    valid_1[290]  <=   0;valid_2[290]  <=   0;dirty_bit_1[290] <= 0;dirty_bit_2[290] <= 0;lru_counter_1[290] <= 0;lru_counter_2[290] <= 0;tag_1[290] <= 0;tag_2[290] <= 0;cache_mem_1[290] <= 0;cache_mem_2[290] <= 0;
    valid_1[291]  <=   0;valid_2[291]  <=   0;dirty_bit_1[291] <= 0;dirty_bit_2[291] <= 0;lru_counter_1[291] <= 0;lru_counter_2[291] <= 0;tag_1[291] <= 0;tag_2[291] <= 0;cache_mem_1[291] <= 0;cache_mem_2[291] <= 0;
    valid_1[292]  <=   0;valid_2[292]  <=   0;dirty_bit_1[292] <= 0;dirty_bit_2[292] <= 0;lru_counter_1[292] <= 0;lru_counter_2[292] <= 0;tag_1[292] <= 0;tag_2[292] <= 0;cache_mem_1[292] <= 0;cache_mem_2[292] <= 0;
    valid_1[293]  <=   0;valid_2[293]  <=   0;dirty_bit_1[293] <= 0;dirty_bit_2[293] <= 0;lru_counter_1[293] <= 0;lru_counter_2[293] <= 0;tag_1[293] <= 0;tag_2[293] <= 0;cache_mem_1[293] <= 0;cache_mem_2[293] <= 0;
    valid_1[294]  <=   0;valid_2[294]  <=   0;dirty_bit_1[294] <= 0;dirty_bit_2[294] <= 0;lru_counter_1[294] <= 0;lru_counter_2[294] <= 0;tag_1[294] <= 0;tag_2[294] <= 0;cache_mem_1[294] <= 0;cache_mem_2[294] <= 0;
    valid_1[295]  <=   0;valid_2[295]  <=   0;dirty_bit_1[295] <= 0;dirty_bit_2[295] <= 0;lru_counter_1[295] <= 0;lru_counter_2[295] <= 0;tag_1[295] <= 0;tag_2[295] <= 0;cache_mem_1[295] <= 0;cache_mem_2[295] <= 0;
    valid_1[296]  <=   0;valid_2[296]  <=   0;dirty_bit_1[296] <= 0;dirty_bit_2[296] <= 0;lru_counter_1[296] <= 0;lru_counter_2[296] <= 0;tag_1[296] <= 0;tag_2[296] <= 0;cache_mem_1[296] <= 0;cache_mem_2[296] <= 0;
    valid_1[297]  <=   0;valid_2[297]  <=   0;dirty_bit_1[297] <= 0;dirty_bit_2[297] <= 0;lru_counter_1[297] <= 0;lru_counter_2[297] <= 0;tag_1[297] <= 0;tag_2[297] <= 0;cache_mem_1[297] <= 0;cache_mem_2[297] <= 0;
    valid_1[298]  <=   0;valid_2[298]  <=   0;dirty_bit_1[298] <= 0;dirty_bit_2[298] <= 0;lru_counter_1[298] <= 0;lru_counter_2[298] <= 0;tag_1[298] <= 0;tag_2[298] <= 0;cache_mem_1[298] <= 0;cache_mem_2[298] <= 0;
    valid_1[299]  <=   0;valid_2[299]  <=   0;dirty_bit_1[299] <= 0;dirty_bit_2[299] <= 0;lru_counter_1[299] <= 0;lru_counter_2[299] <= 0;tag_1[299] <= 0;tag_2[299] <= 0;cache_mem_1[299] <= 0;cache_mem_2[299] <= 0;
    valid_1[300]  <=   0;valid_2[300]  <=   0;dirty_bit_1[300] <= 0;dirty_bit_2[300] <= 0;lru_counter_1[300] <= 0;lru_counter_2[300] <= 0;tag_1[300] <= 0;tag_2[300] <= 0;cache_mem_1[300] <= 0;cache_mem_2[300] <= 0;
    valid_1[301]  <=   0;valid_2[301]  <=   0;dirty_bit_1[301] <= 0;dirty_bit_2[301] <= 0;lru_counter_1[301] <= 0;lru_counter_2[301] <= 0;tag_1[301] <= 0;tag_2[301] <= 0;cache_mem_1[301] <= 0;cache_mem_2[301] <= 0;
    valid_1[302]  <=   0;valid_2[302]  <=   0;dirty_bit_1[302] <= 0;dirty_bit_2[302] <= 0;lru_counter_1[302] <= 0;lru_counter_2[302] <= 0;tag_1[302] <= 0;tag_2[302] <= 0;cache_mem_1[302] <= 0;cache_mem_2[302] <= 0;
    valid_1[303]  <=   0;valid_2[303]  <=   0;dirty_bit_1[303] <= 0;dirty_bit_2[303] <= 0;lru_counter_1[303] <= 0;lru_counter_2[303] <= 0;tag_1[303] <= 0;tag_2[303] <= 0;cache_mem_1[303] <= 0;cache_mem_2[303] <= 0;
    valid_1[304]  <=   0;valid_2[304]  <=   0;dirty_bit_1[304] <= 0;dirty_bit_2[304] <= 0;lru_counter_1[304] <= 0;lru_counter_2[304] <= 0;tag_1[304] <= 0;tag_2[304] <= 0;cache_mem_1[304] <= 0;cache_mem_2[304] <= 0;
    valid_1[305]  <=   0;valid_2[305]  <=   0;dirty_bit_1[305] <= 0;dirty_bit_2[305] <= 0;lru_counter_1[305] <= 0;lru_counter_2[305] <= 0;tag_1[305] <= 0;tag_2[305] <= 0;cache_mem_1[305] <= 0;cache_mem_2[305] <= 0;
    valid_1[306]  <=   0;valid_2[306]  <=   0;dirty_bit_1[306] <= 0;dirty_bit_2[306] <= 0;lru_counter_1[306] <= 0;lru_counter_2[306] <= 0;tag_1[306] <= 0;tag_2[306] <= 0;cache_mem_1[306] <= 0;cache_mem_2[306] <= 0;
    valid_1[307]  <=   0;valid_2[307]  <=   0;dirty_bit_1[307] <= 0;dirty_bit_2[307] <= 0;lru_counter_1[307] <= 0;lru_counter_2[307] <= 0;tag_1[307] <= 0;tag_2[307] <= 0;cache_mem_1[307] <= 0;cache_mem_2[307] <= 0;
    valid_1[308]  <=   0;valid_2[308]  <=   0;dirty_bit_1[308] <= 0;dirty_bit_2[308] <= 0;lru_counter_1[308] <= 0;lru_counter_2[308] <= 0;tag_1[308] <= 0;tag_2[308] <= 0;cache_mem_1[308] <= 0;cache_mem_2[308] <= 0;
    valid_1[309]  <=   0;valid_2[309]  <=   0;dirty_bit_1[309] <= 0;dirty_bit_2[309] <= 0;lru_counter_1[309] <= 0;lru_counter_2[309] <= 0;tag_1[309] <= 0;tag_2[309] <= 0;cache_mem_1[309] <= 0;cache_mem_2[309] <= 0;
    valid_1[310]  <=   0;valid_2[310]  <=   0;dirty_bit_1[310] <= 0;dirty_bit_2[310] <= 0;lru_counter_1[310] <= 0;lru_counter_2[310] <= 0;tag_1[310] <= 0;tag_2[310] <= 0;cache_mem_1[310] <= 0;cache_mem_2[310] <= 0;
    valid_1[311]  <=   0;valid_2[311]  <=   0;dirty_bit_1[311] <= 0;dirty_bit_2[311] <= 0;lru_counter_1[311] <= 0;lru_counter_2[311] <= 0;tag_1[311] <= 0;tag_2[311] <= 0;cache_mem_1[311] <= 0;cache_mem_2[311] <= 0;
    valid_1[312]  <=   0;valid_2[312]  <=   0;dirty_bit_1[312] <= 0;dirty_bit_2[312] <= 0;lru_counter_1[312] <= 0;lru_counter_2[312] <= 0;tag_1[312] <= 0;tag_2[312] <= 0;cache_mem_1[312] <= 0;cache_mem_2[312] <= 0;
    valid_1[313]  <=   0;valid_2[313]  <=   0;dirty_bit_1[313] <= 0;dirty_bit_2[313] <= 0;lru_counter_1[313] <= 0;lru_counter_2[313] <= 0;tag_1[313] <= 0;tag_2[313] <= 0;cache_mem_1[313] <= 0;cache_mem_2[313] <= 0;
    valid_1[314]  <=   0;valid_2[314]  <=   0;dirty_bit_1[314] <= 0;dirty_bit_2[314] <= 0;lru_counter_1[314] <= 0;lru_counter_2[314] <= 0;tag_1[314] <= 0;tag_2[314] <= 0;cache_mem_1[314] <= 0;cache_mem_2[314] <= 0;
    valid_1[315]  <=   0;valid_2[315]  <=   0;dirty_bit_1[315] <= 0;dirty_bit_2[315] <= 0;lru_counter_1[315] <= 0;lru_counter_2[315] <= 0;tag_1[315] <= 0;tag_2[315] <= 0;cache_mem_1[315] <= 0;cache_mem_2[315] <= 0;
    valid_1[316]  <=   0;valid_2[316]  <=   0;dirty_bit_1[316] <= 0;dirty_bit_2[316] <= 0;lru_counter_1[316] <= 0;lru_counter_2[316] <= 0;tag_1[316] <= 0;tag_2[316] <= 0;cache_mem_1[316] <= 0;cache_mem_2[316] <= 0;
    valid_1[317]  <=   0;valid_2[317]  <=   0;dirty_bit_1[317] <= 0;dirty_bit_2[317] <= 0;lru_counter_1[317] <= 0;lru_counter_2[317] <= 0;tag_1[317] <= 0;tag_2[317] <= 0;cache_mem_1[317] <= 0;cache_mem_2[317] <= 0;
    valid_1[318]  <=   0;valid_2[318]  <=   0;dirty_bit_1[318] <= 0;dirty_bit_2[318] <= 0;lru_counter_1[318] <= 0;lru_counter_2[318] <= 0;tag_1[318] <= 0;tag_2[318] <= 0;cache_mem_1[318] <= 0;cache_mem_2[318] <= 0;
    valid_1[319]  <=   0;valid_2[319]  <=   0;dirty_bit_1[319] <= 0;dirty_bit_2[319] <= 0;lru_counter_1[319] <= 0;lru_counter_2[319] <= 0;tag_1[319] <= 0;tag_2[319] <= 0;cache_mem_1[319] <= 0;cache_mem_2[319] <= 0;
    valid_1[320]  <=   0;valid_2[320]  <=   0;dirty_bit_1[320] <= 0;dirty_bit_2[320] <= 0;lru_counter_1[320] <= 0;lru_counter_2[320] <= 0;tag_1[320] <= 0;tag_2[320] <= 0;cache_mem_1[320] <= 0;cache_mem_2[320] <= 0;
    valid_1[321]  <=   0;valid_2[321]  <=   0;dirty_bit_1[321] <= 0;dirty_bit_2[321] <= 0;lru_counter_1[321] <= 0;lru_counter_2[321] <= 0;tag_1[321] <= 0;tag_2[321] <= 0;cache_mem_1[321] <= 0;cache_mem_2[321] <= 0;
    valid_1[322]  <=   0;valid_2[322]  <=   0;dirty_bit_1[322] <= 0;dirty_bit_2[322] <= 0;lru_counter_1[322] <= 0;lru_counter_2[322] <= 0;tag_1[322] <= 0;tag_2[322] <= 0;cache_mem_1[322] <= 0;cache_mem_2[322] <= 0;
    valid_1[323]  <=   0;valid_2[323]  <=   0;dirty_bit_1[323] <= 0;dirty_bit_2[323] <= 0;lru_counter_1[323] <= 0;lru_counter_2[323] <= 0;tag_1[323] <= 0;tag_2[323] <= 0;cache_mem_1[323] <= 0;cache_mem_2[323] <= 0;
    valid_1[324]  <=   0;valid_2[324]  <=   0;dirty_bit_1[324] <= 0;dirty_bit_2[324] <= 0;lru_counter_1[324] <= 0;lru_counter_2[324] <= 0;tag_1[324] <= 0;tag_2[324] <= 0;cache_mem_1[324] <= 0;cache_mem_2[324] <= 0;
    valid_1[325]  <=   0;valid_2[325]  <=   0;dirty_bit_1[325] <= 0;dirty_bit_2[325] <= 0;lru_counter_1[325] <= 0;lru_counter_2[325] <= 0;tag_1[325] <= 0;tag_2[325] <= 0;cache_mem_1[325] <= 0;cache_mem_2[325] <= 0;
    valid_1[326]  <=   0;valid_2[326]  <=   0;dirty_bit_1[326] <= 0;dirty_bit_2[326] <= 0;lru_counter_1[326] <= 0;lru_counter_2[326] <= 0;tag_1[326] <= 0;tag_2[326] <= 0;cache_mem_1[326] <= 0;cache_mem_2[326] <= 0;
    valid_1[327]  <=   0;valid_2[327]  <=   0;dirty_bit_1[327] <= 0;dirty_bit_2[327] <= 0;lru_counter_1[327] <= 0;lru_counter_2[327] <= 0;tag_1[327] <= 0;tag_2[327] <= 0;cache_mem_1[327] <= 0;cache_mem_2[327] <= 0;
    valid_1[328]  <=   0;valid_2[328]  <=   0;dirty_bit_1[328] <= 0;dirty_bit_2[328] <= 0;lru_counter_1[328] <= 0;lru_counter_2[328] <= 0;tag_1[328] <= 0;tag_2[328] <= 0;cache_mem_1[328] <= 0;cache_mem_2[328] <= 0;
    valid_1[329]  <=   0;valid_2[329]  <=   0;dirty_bit_1[329] <= 0;dirty_bit_2[329] <= 0;lru_counter_1[329] <= 0;lru_counter_2[329] <= 0;tag_1[329] <= 0;tag_2[329] <= 0;cache_mem_1[329] <= 0;cache_mem_2[329] <= 0;
    valid_1[330]  <=   0;valid_2[330]  <=   0;dirty_bit_1[330] <= 0;dirty_bit_2[330] <= 0;lru_counter_1[330] <= 0;lru_counter_2[330] <= 0;tag_1[330] <= 0;tag_2[330] <= 0;cache_mem_1[330] <= 0;cache_mem_2[330] <= 0;
    valid_1[331]  <=   0;valid_2[331]  <=   0;dirty_bit_1[331] <= 0;dirty_bit_2[331] <= 0;lru_counter_1[331] <= 0;lru_counter_2[331] <= 0;tag_1[331] <= 0;tag_2[331] <= 0;cache_mem_1[331] <= 0;cache_mem_2[331] <= 0;
    valid_1[332]  <=   0;valid_2[332]  <=   0;dirty_bit_1[332] <= 0;dirty_bit_2[332] <= 0;lru_counter_1[332] <= 0;lru_counter_2[332] <= 0;tag_1[332] <= 0;tag_2[332] <= 0;cache_mem_1[332] <= 0;cache_mem_2[332] <= 0;
    valid_1[333]  <=   0;valid_2[333]  <=   0;dirty_bit_1[333] <= 0;dirty_bit_2[333] <= 0;lru_counter_1[333] <= 0;lru_counter_2[333] <= 0;tag_1[333] <= 0;tag_2[333] <= 0;cache_mem_1[333] <= 0;cache_mem_2[333] <= 0;
    valid_1[334]  <=   0;valid_2[334]  <=   0;dirty_bit_1[334] <= 0;dirty_bit_2[334] <= 0;lru_counter_1[334] <= 0;lru_counter_2[334] <= 0;tag_1[334] <= 0;tag_2[334] <= 0;cache_mem_1[334] <= 0;cache_mem_2[334] <= 0;
    valid_1[335]  <=   0;valid_2[335]  <=   0;dirty_bit_1[335] <= 0;dirty_bit_2[335] <= 0;lru_counter_1[335] <= 0;lru_counter_2[335] <= 0;tag_1[335] <= 0;tag_2[335] <= 0;cache_mem_1[335] <= 0;cache_mem_2[335] <= 0;
    valid_1[336]  <=   0;valid_2[336]  <=   0;dirty_bit_1[336] <= 0;dirty_bit_2[336] <= 0;lru_counter_1[336] <= 0;lru_counter_2[336] <= 0;tag_1[336] <= 0;tag_2[336] <= 0;cache_mem_1[336] <= 0;cache_mem_2[336] <= 0;
    valid_1[337]  <=   0;valid_2[337]  <=   0;dirty_bit_1[337] <= 0;dirty_bit_2[337] <= 0;lru_counter_1[337] <= 0;lru_counter_2[337] <= 0;tag_1[337] <= 0;tag_2[337] <= 0;cache_mem_1[337] <= 0;cache_mem_2[337] <= 0;
    valid_1[338]  <=   0;valid_2[338]  <=   0;dirty_bit_1[338] <= 0;dirty_bit_2[338] <= 0;lru_counter_1[338] <= 0;lru_counter_2[338] <= 0;tag_1[338] <= 0;tag_2[338] <= 0;cache_mem_1[338] <= 0;cache_mem_2[338] <= 0;
    valid_1[339]  <=   0;valid_2[339]  <=   0;dirty_bit_1[339] <= 0;dirty_bit_2[339] <= 0;lru_counter_1[339] <= 0;lru_counter_2[339] <= 0;tag_1[339] <= 0;tag_2[339] <= 0;cache_mem_1[339] <= 0;cache_mem_2[339] <= 0;
    valid_1[340]  <=   0;valid_2[340]  <=   0;dirty_bit_1[340] <= 0;dirty_bit_2[340] <= 0;lru_counter_1[340] <= 0;lru_counter_2[340] <= 0;tag_1[340] <= 0;tag_2[340] <= 0;cache_mem_1[340] <= 0;cache_mem_2[340] <= 0;
    valid_1[341]  <=   0;valid_2[341]  <=   0;dirty_bit_1[341] <= 0;dirty_bit_2[341] <= 0;lru_counter_1[341] <= 0;lru_counter_2[341] <= 0;tag_1[341] <= 0;tag_2[341] <= 0;cache_mem_1[341] <= 0;cache_mem_2[341] <= 0;
    valid_1[342]  <=   0;valid_2[342]  <=   0;dirty_bit_1[342] <= 0;dirty_bit_2[342] <= 0;lru_counter_1[342] <= 0;lru_counter_2[342] <= 0;tag_1[342] <= 0;tag_2[342] <= 0;cache_mem_1[342] <= 0;cache_mem_2[342] <= 0;
    valid_1[343]  <=   0;valid_2[343]  <=   0;dirty_bit_1[343] <= 0;dirty_bit_2[343] <= 0;lru_counter_1[343] <= 0;lru_counter_2[343] <= 0;tag_1[343] <= 0;tag_2[343] <= 0;cache_mem_1[343] <= 0;cache_mem_2[343] <= 0;
    valid_1[344]  <=   0;valid_2[344]  <=   0;dirty_bit_1[344] <= 0;dirty_bit_2[344] <= 0;lru_counter_1[344] <= 0;lru_counter_2[344] <= 0;tag_1[344] <= 0;tag_2[344] <= 0;cache_mem_1[344] <= 0;cache_mem_2[344] <= 0;
    valid_1[345]  <=   0;valid_2[345]  <=   0;dirty_bit_1[345] <= 0;dirty_bit_2[345] <= 0;lru_counter_1[345] <= 0;lru_counter_2[345] <= 0;tag_1[345] <= 0;tag_2[345] <= 0;cache_mem_1[345] <= 0;cache_mem_2[345] <= 0;
    valid_1[346]  <=   0;valid_2[346]  <=   0;dirty_bit_1[346] <= 0;dirty_bit_2[346] <= 0;lru_counter_1[346] <= 0;lru_counter_2[346] <= 0;tag_1[346] <= 0;tag_2[346] <= 0;cache_mem_1[346] <= 0;cache_mem_2[346] <= 0;
    valid_1[347]  <=   0;valid_2[347]  <=   0;dirty_bit_1[347] <= 0;dirty_bit_2[347] <= 0;lru_counter_1[347] <= 0;lru_counter_2[347] <= 0;tag_1[347] <= 0;tag_2[347] <= 0;cache_mem_1[347] <= 0;cache_mem_2[347] <= 0;
    valid_1[348]  <=   0;valid_2[348]  <=   0;dirty_bit_1[348] <= 0;dirty_bit_2[348] <= 0;lru_counter_1[348] <= 0;lru_counter_2[348] <= 0;tag_1[348] <= 0;tag_2[348] <= 0;cache_mem_1[348] <= 0;cache_mem_2[348] <= 0;
    valid_1[349]  <=   0;valid_2[349]  <=   0;dirty_bit_1[349] <= 0;dirty_bit_2[349] <= 0;lru_counter_1[349] <= 0;lru_counter_2[349] <= 0;tag_1[349] <= 0;tag_2[349] <= 0;cache_mem_1[349] <= 0;cache_mem_2[349] <= 0;
    valid_1[350]  <=   0;valid_2[350]  <=   0;dirty_bit_1[350] <= 0;dirty_bit_2[350] <= 0;lru_counter_1[350] <= 0;lru_counter_2[350] <= 0;tag_1[350] <= 0;tag_2[350] <= 0;cache_mem_1[350] <= 0;cache_mem_2[350] <= 0;
    valid_1[351]  <=   0;valid_2[351]  <=   0;dirty_bit_1[351] <= 0;dirty_bit_2[351] <= 0;lru_counter_1[351] <= 0;lru_counter_2[351] <= 0;tag_1[351] <= 0;tag_2[351] <= 0;cache_mem_1[351] <= 0;cache_mem_2[351] <= 0;
    valid_1[352]  <=   0;valid_2[352]  <=   0;dirty_bit_1[352] <= 0;dirty_bit_2[352] <= 0;lru_counter_1[352] <= 0;lru_counter_2[352] <= 0;tag_1[352] <= 0;tag_2[352] <= 0;cache_mem_1[352] <= 0;cache_mem_2[352] <= 0;
    valid_1[353]  <=   0;valid_2[353]  <=   0;dirty_bit_1[353] <= 0;dirty_bit_2[353] <= 0;lru_counter_1[353] <= 0;lru_counter_2[353] <= 0;tag_1[353] <= 0;tag_2[353] <= 0;cache_mem_1[353] <= 0;cache_mem_2[353] <= 0;
    valid_1[354]  <=   0;valid_2[354]  <=   0;dirty_bit_1[354] <= 0;dirty_bit_2[354] <= 0;lru_counter_1[354] <= 0;lru_counter_2[354] <= 0;tag_1[354] <= 0;tag_2[354] <= 0;cache_mem_1[354] <= 0;cache_mem_2[354] <= 0;
    valid_1[355]  <=   0;valid_2[355]  <=   0;dirty_bit_1[355] <= 0;dirty_bit_2[355] <= 0;lru_counter_1[355] <= 0;lru_counter_2[355] <= 0;tag_1[355] <= 0;tag_2[355] <= 0;cache_mem_1[355] <= 0;cache_mem_2[355] <= 0;
    valid_1[356]  <=   0;valid_2[356]  <=   0;dirty_bit_1[356] <= 0;dirty_bit_2[356] <= 0;lru_counter_1[356] <= 0;lru_counter_2[356] <= 0;tag_1[356] <= 0;tag_2[356] <= 0;cache_mem_1[356] <= 0;cache_mem_2[356] <= 0;
    valid_1[357]  <=   0;valid_2[357]  <=   0;dirty_bit_1[357] <= 0;dirty_bit_2[357] <= 0;lru_counter_1[357] <= 0;lru_counter_2[357] <= 0;tag_1[357] <= 0;tag_2[357] <= 0;cache_mem_1[357] <= 0;cache_mem_2[357] <= 0;
    valid_1[358]  <=   0;valid_2[358]  <=   0;dirty_bit_1[358] <= 0;dirty_bit_2[358] <= 0;lru_counter_1[358] <= 0;lru_counter_2[358] <= 0;tag_1[358] <= 0;tag_2[358] <= 0;cache_mem_1[358] <= 0;cache_mem_2[358] <= 0;
    valid_1[359]  <=   0;valid_2[359]  <=   0;dirty_bit_1[359] <= 0;dirty_bit_2[359] <= 0;lru_counter_1[359] <= 0;lru_counter_2[359] <= 0;tag_1[359] <= 0;tag_2[359] <= 0;cache_mem_1[359] <= 0;cache_mem_2[359] <= 0;
    valid_1[360]  <=   0;valid_2[360]  <=   0;dirty_bit_1[360] <= 0;dirty_bit_2[360] <= 0;lru_counter_1[360] <= 0;lru_counter_2[360] <= 0;tag_1[360] <= 0;tag_2[360] <= 0;cache_mem_1[360] <= 0;cache_mem_2[360] <= 0;
    valid_1[361]  <=   0;valid_2[361]  <=   0;dirty_bit_1[361] <= 0;dirty_bit_2[361] <= 0;lru_counter_1[361] <= 0;lru_counter_2[361] <= 0;tag_1[361] <= 0;tag_2[361] <= 0;cache_mem_1[361] <= 0;cache_mem_2[361] <= 0;
    valid_1[362]  <=   0;valid_2[362]  <=   0;dirty_bit_1[362] <= 0;dirty_bit_2[362] <= 0;lru_counter_1[362] <= 0;lru_counter_2[362] <= 0;tag_1[362] <= 0;tag_2[362] <= 0;cache_mem_1[362] <= 0;cache_mem_2[362] <= 0;
    valid_1[363]  <=   0;valid_2[363]  <=   0;dirty_bit_1[363] <= 0;dirty_bit_2[363] <= 0;lru_counter_1[363] <= 0;lru_counter_2[363] <= 0;tag_1[363] <= 0;tag_2[363] <= 0;cache_mem_1[363] <= 0;cache_mem_2[363] <= 0;
    valid_1[364]  <=   0;valid_2[364]  <=   0;dirty_bit_1[364] <= 0;dirty_bit_2[364] <= 0;lru_counter_1[364] <= 0;lru_counter_2[364] <= 0;tag_1[364] <= 0;tag_2[364] <= 0;cache_mem_1[364] <= 0;cache_mem_2[364] <= 0;
    valid_1[365]  <=   0;valid_2[365]  <=   0;dirty_bit_1[365] <= 0;dirty_bit_2[365] <= 0;lru_counter_1[365] <= 0;lru_counter_2[365] <= 0;tag_1[365] <= 0;tag_2[365] <= 0;cache_mem_1[365] <= 0;cache_mem_2[365] <= 0;
    valid_1[366]  <=   0;valid_2[366]  <=   0;dirty_bit_1[366] <= 0;dirty_bit_2[366] <= 0;lru_counter_1[366] <= 0;lru_counter_2[366] <= 0;tag_1[366] <= 0;tag_2[366] <= 0;cache_mem_1[366] <= 0;cache_mem_2[366] <= 0;
    valid_1[367]  <=   0;valid_2[367]  <=   0;dirty_bit_1[367] <= 0;dirty_bit_2[367] <= 0;lru_counter_1[367] <= 0;lru_counter_2[367] <= 0;tag_1[367] <= 0;tag_2[367] <= 0;cache_mem_1[367] <= 0;cache_mem_2[367] <= 0;
    valid_1[368]  <=   0;valid_2[368]  <=   0;dirty_bit_1[368] <= 0;dirty_bit_2[368] <= 0;lru_counter_1[368] <= 0;lru_counter_2[368] <= 0;tag_1[368] <= 0;tag_2[368] <= 0;cache_mem_1[368] <= 0;cache_mem_2[368] <= 0;
    valid_1[369]  <=   0;valid_2[369]  <=   0;dirty_bit_1[369] <= 0;dirty_bit_2[369] <= 0;lru_counter_1[369] <= 0;lru_counter_2[369] <= 0;tag_1[369] <= 0;tag_2[369] <= 0;cache_mem_1[369] <= 0;cache_mem_2[369] <= 0;
    valid_1[370]  <=   0;valid_2[370]  <=   0;dirty_bit_1[370] <= 0;dirty_bit_2[370] <= 0;lru_counter_1[370] <= 0;lru_counter_2[370] <= 0;tag_1[370] <= 0;tag_2[370] <= 0;cache_mem_1[370] <= 0;cache_mem_2[370] <= 0;
    valid_1[371]  <=   0;valid_2[371]  <=   0;dirty_bit_1[371] <= 0;dirty_bit_2[371] <= 0;lru_counter_1[371] <= 0;lru_counter_2[371] <= 0;tag_1[371] <= 0;tag_2[371] <= 0;cache_mem_1[371] <= 0;cache_mem_2[371] <= 0;
    valid_1[372]  <=   0;valid_2[372]  <=   0;dirty_bit_1[372] <= 0;dirty_bit_2[372] <= 0;lru_counter_1[372] <= 0;lru_counter_2[372] <= 0;tag_1[372] <= 0;tag_2[372] <= 0;cache_mem_1[372] <= 0;cache_mem_2[372] <= 0;
    valid_1[373]  <=   0;valid_2[373]  <=   0;dirty_bit_1[373] <= 0;dirty_bit_2[373] <= 0;lru_counter_1[373] <= 0;lru_counter_2[373] <= 0;tag_1[373] <= 0;tag_2[373] <= 0;cache_mem_1[373] <= 0;cache_mem_2[373] <= 0;
    valid_1[374]  <=   0;valid_2[374]  <=   0;dirty_bit_1[374] <= 0;dirty_bit_2[374] <= 0;lru_counter_1[374] <= 0;lru_counter_2[374] <= 0;tag_1[374] <= 0;tag_2[374] <= 0;cache_mem_1[374] <= 0;cache_mem_2[374] <= 0;
    valid_1[375]  <=   0;valid_2[375]  <=   0;dirty_bit_1[375] <= 0;dirty_bit_2[375] <= 0;lru_counter_1[375] <= 0;lru_counter_2[375] <= 0;tag_1[375] <= 0;tag_2[375] <= 0;cache_mem_1[375] <= 0;cache_mem_2[375] <= 0;
    valid_1[376]  <=   0;valid_2[376]  <=   0;dirty_bit_1[376] <= 0;dirty_bit_2[376] <= 0;lru_counter_1[376] <= 0;lru_counter_2[376] <= 0;tag_1[376] <= 0;tag_2[376] <= 0;cache_mem_1[376] <= 0;cache_mem_2[376] <= 0;
    valid_1[377]  <=   0;valid_2[377]  <=   0;dirty_bit_1[377] <= 0;dirty_bit_2[377] <= 0;lru_counter_1[377] <= 0;lru_counter_2[377] <= 0;tag_1[377] <= 0;tag_2[377] <= 0;cache_mem_1[377] <= 0;cache_mem_2[377] <= 0;
    valid_1[378]  <=   0;valid_2[378]  <=   0;dirty_bit_1[378] <= 0;dirty_bit_2[378] <= 0;lru_counter_1[378] <= 0;lru_counter_2[378] <= 0;tag_1[378] <= 0;tag_2[378] <= 0;cache_mem_1[378] <= 0;cache_mem_2[378] <= 0;
    valid_1[379]  <=   0;valid_2[379]  <=   0;dirty_bit_1[379] <= 0;dirty_bit_2[379] <= 0;lru_counter_1[379] <= 0;lru_counter_2[379] <= 0;tag_1[379] <= 0;tag_2[379] <= 0;cache_mem_1[379] <= 0;cache_mem_2[379] <= 0;
    valid_1[380]  <=   0;valid_2[380]  <=   0;dirty_bit_1[380] <= 0;dirty_bit_2[380] <= 0;lru_counter_1[380] <= 0;lru_counter_2[380] <= 0;tag_1[380] <= 0;tag_2[380] <= 0;cache_mem_1[380] <= 0;cache_mem_2[380] <= 0;
    valid_1[381]  <=   0;valid_2[381]  <=   0;dirty_bit_1[381] <= 0;dirty_bit_2[381] <= 0;lru_counter_1[381] <= 0;lru_counter_2[381] <= 0;tag_1[381] <= 0;tag_2[381] <= 0;cache_mem_1[381] <= 0;cache_mem_2[381] <= 0;
    valid_1[382]  <=   0;valid_2[382]  <=   0;dirty_bit_1[382] <= 0;dirty_bit_2[382] <= 0;lru_counter_1[382] <= 0;lru_counter_2[382] <= 0;tag_1[382] <= 0;tag_2[382] <= 0;cache_mem_1[382] <= 0;cache_mem_2[382] <= 0;
    valid_1[383]  <=   0;valid_2[383]  <=   0;dirty_bit_1[383] <= 0;dirty_bit_2[383] <= 0;lru_counter_1[383] <= 0;lru_counter_2[383] <= 0;tag_1[383] <= 0;tag_2[383] <= 0;cache_mem_1[383] <= 0;cache_mem_2[383] <= 0;
    valid_1[384]  <=   0;valid_2[384]  <=   0;dirty_bit_1[384] <= 0;dirty_bit_2[384] <= 0;lru_counter_1[384] <= 0;lru_counter_2[384] <= 0;tag_1[384] <= 0;tag_2[384] <= 0;cache_mem_1[384] <= 0;cache_mem_2[384] <= 0;
    valid_1[385]  <=   0;valid_2[385]  <=   0;dirty_bit_1[385] <= 0;dirty_bit_2[385] <= 0;lru_counter_1[385] <= 0;lru_counter_2[385] <= 0;tag_1[385] <= 0;tag_2[385] <= 0;cache_mem_1[385] <= 0;cache_mem_2[385] <= 0;
    valid_1[386]  <=   0;valid_2[386]  <=   0;dirty_bit_1[386] <= 0;dirty_bit_2[386] <= 0;lru_counter_1[386] <= 0;lru_counter_2[386] <= 0;tag_1[386] <= 0;tag_2[386] <= 0;cache_mem_1[386] <= 0;cache_mem_2[386] <= 0;
    valid_1[387]  <=   0;valid_2[387]  <=   0;dirty_bit_1[387] <= 0;dirty_bit_2[387] <= 0;lru_counter_1[387] <= 0;lru_counter_2[387] <= 0;tag_1[387] <= 0;tag_2[387] <= 0;cache_mem_1[387] <= 0;cache_mem_2[387] <= 0;
    valid_1[388]  <=   0;valid_2[388]  <=   0;dirty_bit_1[388] <= 0;dirty_bit_2[388] <= 0;lru_counter_1[388] <= 0;lru_counter_2[388] <= 0;tag_1[388] <= 0;tag_2[388] <= 0;cache_mem_1[388] <= 0;cache_mem_2[388] <= 0;
    valid_1[389]  <=   0;valid_2[389]  <=   0;dirty_bit_1[389] <= 0;dirty_bit_2[389] <= 0;lru_counter_1[389] <= 0;lru_counter_2[389] <= 0;tag_1[389] <= 0;tag_2[389] <= 0;cache_mem_1[389] <= 0;cache_mem_2[389] <= 0;
    valid_1[390]  <=   0;valid_2[390]  <=   0;dirty_bit_1[390] <= 0;dirty_bit_2[390] <= 0;lru_counter_1[390] <= 0;lru_counter_2[390] <= 0;tag_1[390] <= 0;tag_2[390] <= 0;cache_mem_1[390] <= 0;cache_mem_2[390] <= 0;
    valid_1[391]  <=   0;valid_2[391]  <=   0;dirty_bit_1[391] <= 0;dirty_bit_2[391] <= 0;lru_counter_1[391] <= 0;lru_counter_2[391] <= 0;tag_1[391] <= 0;tag_2[391] <= 0;cache_mem_1[391] <= 0;cache_mem_2[391] <= 0;
    valid_1[392]  <=   0;valid_2[392]  <=   0;dirty_bit_1[392] <= 0;dirty_bit_2[392] <= 0;lru_counter_1[392] <= 0;lru_counter_2[392] <= 0;tag_1[392] <= 0;tag_2[392] <= 0;cache_mem_1[392] <= 0;cache_mem_2[392] <= 0;
    valid_1[393]  <=   0;valid_2[393]  <=   0;dirty_bit_1[393] <= 0;dirty_bit_2[393] <= 0;lru_counter_1[393] <= 0;lru_counter_2[393] <= 0;tag_1[393] <= 0;tag_2[393] <= 0;cache_mem_1[393] <= 0;cache_mem_2[393] <= 0;
    valid_1[394]  <=   0;valid_2[394]  <=   0;dirty_bit_1[394] <= 0;dirty_bit_2[394] <= 0;lru_counter_1[394] <= 0;lru_counter_2[394] <= 0;tag_1[394] <= 0;tag_2[394] <= 0;cache_mem_1[394] <= 0;cache_mem_2[394] <= 0;
    valid_1[395]  <=   0;valid_2[395]  <=   0;dirty_bit_1[395] <= 0;dirty_bit_2[395] <= 0;lru_counter_1[395] <= 0;lru_counter_2[395] <= 0;tag_1[395] <= 0;tag_2[395] <= 0;cache_mem_1[395] <= 0;cache_mem_2[395] <= 0;
    valid_1[396]  <=   0;valid_2[396]  <=   0;dirty_bit_1[396] <= 0;dirty_bit_2[396] <= 0;lru_counter_1[396] <= 0;lru_counter_2[396] <= 0;tag_1[396] <= 0;tag_2[396] <= 0;cache_mem_1[396] <= 0;cache_mem_2[396] <= 0;
    valid_1[397]  <=   0;valid_2[397]  <=   0;dirty_bit_1[397] <= 0;dirty_bit_2[397] <= 0;lru_counter_1[397] <= 0;lru_counter_2[397] <= 0;tag_1[397] <= 0;tag_2[397] <= 0;cache_mem_1[397] <= 0;cache_mem_2[397] <= 0;
    valid_1[398]  <=   0;valid_2[398]  <=   0;dirty_bit_1[398] <= 0;dirty_bit_2[398] <= 0;lru_counter_1[398] <= 0;lru_counter_2[398] <= 0;tag_1[398] <= 0;tag_2[398] <= 0;cache_mem_1[398] <= 0;cache_mem_2[398] <= 0;
    valid_1[399]  <=   0;valid_2[399]  <=   0;dirty_bit_1[399] <= 0;dirty_bit_2[399] <= 0;lru_counter_1[399] <= 0;lru_counter_2[399] <= 0;tag_1[399] <= 0;tag_2[399] <= 0;cache_mem_1[399] <= 0;cache_mem_2[399] <= 0;
    valid_1[400]  <=   0;valid_2[400]  <=   0;dirty_bit_1[400] <= 0;dirty_bit_2[400] <= 0;lru_counter_1[400] <= 0;lru_counter_2[400] <= 0;tag_1[400] <= 0;tag_2[400] <= 0;cache_mem_1[400] <= 0;cache_mem_2[400] <= 0;
    valid_1[401]  <=   0;valid_2[401]  <=   0;dirty_bit_1[401] <= 0;dirty_bit_2[401] <= 0;lru_counter_1[401] <= 0;lru_counter_2[401] <= 0;tag_1[401] <= 0;tag_2[401] <= 0;cache_mem_1[401] <= 0;cache_mem_2[401] <= 0;
    valid_1[402]  <=   0;valid_2[402]  <=   0;dirty_bit_1[402] <= 0;dirty_bit_2[402] <= 0;lru_counter_1[402] <= 0;lru_counter_2[402] <= 0;tag_1[402] <= 0;tag_2[402] <= 0;cache_mem_1[402] <= 0;cache_mem_2[402] <= 0;
    valid_1[403]  <=   0;valid_2[403]  <=   0;dirty_bit_1[403] <= 0;dirty_bit_2[403] <= 0;lru_counter_1[403] <= 0;lru_counter_2[403] <= 0;tag_1[403] <= 0;tag_2[403] <= 0;cache_mem_1[403] <= 0;cache_mem_2[403] <= 0;
    valid_1[404]  <=   0;valid_2[404]  <=   0;dirty_bit_1[404] <= 0;dirty_bit_2[404] <= 0;lru_counter_1[404] <= 0;lru_counter_2[404] <= 0;tag_1[404] <= 0;tag_2[404] <= 0;cache_mem_1[404] <= 0;cache_mem_2[404] <= 0;
    valid_1[405]  <=   0;valid_2[405]  <=   0;dirty_bit_1[405] <= 0;dirty_bit_2[405] <= 0;lru_counter_1[405] <= 0;lru_counter_2[405] <= 0;tag_1[405] <= 0;tag_2[405] <= 0;cache_mem_1[405] <= 0;cache_mem_2[405] <= 0;
    valid_1[406]  <=   0;valid_2[406]  <=   0;dirty_bit_1[406] <= 0;dirty_bit_2[406] <= 0;lru_counter_1[406] <= 0;lru_counter_2[406] <= 0;tag_1[406] <= 0;tag_2[406] <= 0;cache_mem_1[406] <= 0;cache_mem_2[406] <= 0;
    valid_1[407]  <=   0;valid_2[407]  <=   0;dirty_bit_1[407] <= 0;dirty_bit_2[407] <= 0;lru_counter_1[407] <= 0;lru_counter_2[407] <= 0;tag_1[407] <= 0;tag_2[407] <= 0;cache_mem_1[407] <= 0;cache_mem_2[407] <= 0;
    valid_1[408]  <=   0;valid_2[408]  <=   0;dirty_bit_1[408] <= 0;dirty_bit_2[408] <= 0;lru_counter_1[408] <= 0;lru_counter_2[408] <= 0;tag_1[408] <= 0;tag_2[408] <= 0;cache_mem_1[408] <= 0;cache_mem_2[408] <= 0;
    valid_1[409]  <=   0;valid_2[409]  <=   0;dirty_bit_1[409] <= 0;dirty_bit_2[409] <= 0;lru_counter_1[409] <= 0;lru_counter_2[409] <= 0;tag_1[409] <= 0;tag_2[409] <= 0;cache_mem_1[409] <= 0;cache_mem_2[409] <= 0;
    valid_1[410]  <=   0;valid_2[410]  <=   0;dirty_bit_1[410] <= 0;dirty_bit_2[410] <= 0;lru_counter_1[410] <= 0;lru_counter_2[410] <= 0;tag_1[410] <= 0;tag_2[410] <= 0;cache_mem_1[410] <= 0;cache_mem_2[410] <= 0;
    valid_1[411]  <=   0;valid_2[411]  <=   0;dirty_bit_1[411] <= 0;dirty_bit_2[411] <= 0;lru_counter_1[411] <= 0;lru_counter_2[411] <= 0;tag_1[411] <= 0;tag_2[411] <= 0;cache_mem_1[411] <= 0;cache_mem_2[411] <= 0;
    valid_1[412]  <=   0;valid_2[412]  <=   0;dirty_bit_1[412] <= 0;dirty_bit_2[412] <= 0;lru_counter_1[412] <= 0;lru_counter_2[412] <= 0;tag_1[412] <= 0;tag_2[412] <= 0;cache_mem_1[412] <= 0;cache_mem_2[412] <= 0;
    valid_1[413]  <=   0;valid_2[413]  <=   0;dirty_bit_1[413] <= 0;dirty_bit_2[413] <= 0;lru_counter_1[413] <= 0;lru_counter_2[413] <= 0;tag_1[413] <= 0;tag_2[413] <= 0;cache_mem_1[413] <= 0;cache_mem_2[413] <= 0;
    valid_1[414]  <=   0;valid_2[414]  <=   0;dirty_bit_1[414] <= 0;dirty_bit_2[414] <= 0;lru_counter_1[414] <= 0;lru_counter_2[414] <= 0;tag_1[414] <= 0;tag_2[414] <= 0;cache_mem_1[414] <= 0;cache_mem_2[414] <= 0;
    valid_1[415]  <=   0;valid_2[415]  <=   0;dirty_bit_1[415] <= 0;dirty_bit_2[415] <= 0;lru_counter_1[415] <= 0;lru_counter_2[415] <= 0;tag_1[415] <= 0;tag_2[415] <= 0;cache_mem_1[415] <= 0;cache_mem_2[415] <= 0;
    valid_1[416]  <=   0;valid_2[416]  <=   0;dirty_bit_1[416] <= 0;dirty_bit_2[416] <= 0;lru_counter_1[416] <= 0;lru_counter_2[416] <= 0;tag_1[416] <= 0;tag_2[416] <= 0;cache_mem_1[416] <= 0;cache_mem_2[416] <= 0;
    valid_1[417]  <=   0;valid_2[417]  <=   0;dirty_bit_1[417] <= 0;dirty_bit_2[417] <= 0;lru_counter_1[417] <= 0;lru_counter_2[417] <= 0;tag_1[417] <= 0;tag_2[417] <= 0;cache_mem_1[417] <= 0;cache_mem_2[417] <= 0;
    valid_1[418]  <=   0;valid_2[418]  <=   0;dirty_bit_1[418] <= 0;dirty_bit_2[418] <= 0;lru_counter_1[418] <= 0;lru_counter_2[418] <= 0;tag_1[418] <= 0;tag_2[418] <= 0;cache_mem_1[418] <= 0;cache_mem_2[418] <= 0;
    valid_1[419]  <=   0;valid_2[419]  <=   0;dirty_bit_1[419] <= 0;dirty_bit_2[419] <= 0;lru_counter_1[419] <= 0;lru_counter_2[419] <= 0;tag_1[419] <= 0;tag_2[419] <= 0;cache_mem_1[419] <= 0;cache_mem_2[419] <= 0;
    valid_1[420]  <=   0;valid_2[420]  <=   0;dirty_bit_1[420] <= 0;dirty_bit_2[420] <= 0;lru_counter_1[420] <= 0;lru_counter_2[420] <= 0;tag_1[420] <= 0;tag_2[420] <= 0;cache_mem_1[420] <= 0;cache_mem_2[420] <= 0;
    valid_1[421]  <=   0;valid_2[421]  <=   0;dirty_bit_1[421] <= 0;dirty_bit_2[421] <= 0;lru_counter_1[421] <= 0;lru_counter_2[421] <= 0;tag_1[421] <= 0;tag_2[421] <= 0;cache_mem_1[421] <= 0;cache_mem_2[421] <= 0;
    valid_1[422]  <=   0;valid_2[422]  <=   0;dirty_bit_1[422] <= 0;dirty_bit_2[422] <= 0;lru_counter_1[422] <= 0;lru_counter_2[422] <= 0;tag_1[422] <= 0;tag_2[422] <= 0;cache_mem_1[422] <= 0;cache_mem_2[422] <= 0;
    valid_1[423]  <=   0;valid_2[423]  <=   0;dirty_bit_1[423] <= 0;dirty_bit_2[423] <= 0;lru_counter_1[423] <= 0;lru_counter_2[423] <= 0;tag_1[423] <= 0;tag_2[423] <= 0;cache_mem_1[423] <= 0;cache_mem_2[423] <= 0;
    valid_1[424]  <=   0;valid_2[424]  <=   0;dirty_bit_1[424] <= 0;dirty_bit_2[424] <= 0;lru_counter_1[424] <= 0;lru_counter_2[424] <= 0;tag_1[424] <= 0;tag_2[424] <= 0;cache_mem_1[424] <= 0;cache_mem_2[424] <= 0;
    valid_1[425]  <=   0;valid_2[425]  <=   0;dirty_bit_1[425] <= 0;dirty_bit_2[425] <= 0;lru_counter_1[425] <= 0;lru_counter_2[425] <= 0;tag_1[425] <= 0;tag_2[425] <= 0;cache_mem_1[425] <= 0;cache_mem_2[425] <= 0;
    valid_1[426]  <=   0;valid_2[426]  <=   0;dirty_bit_1[426] <= 0;dirty_bit_2[426] <= 0;lru_counter_1[426] <= 0;lru_counter_2[426] <= 0;tag_1[426] <= 0;tag_2[426] <= 0;cache_mem_1[426] <= 0;cache_mem_2[426] <= 0;
    valid_1[427]  <=   0;valid_2[427]  <=   0;dirty_bit_1[427] <= 0;dirty_bit_2[427] <= 0;lru_counter_1[427] <= 0;lru_counter_2[427] <= 0;tag_1[427] <= 0;tag_2[427] <= 0;cache_mem_1[427] <= 0;cache_mem_2[427] <= 0;
    valid_1[428]  <=   0;valid_2[428]  <=   0;dirty_bit_1[428] <= 0;dirty_bit_2[428] <= 0;lru_counter_1[428] <= 0;lru_counter_2[428] <= 0;tag_1[428] <= 0;tag_2[428] <= 0;cache_mem_1[428] <= 0;cache_mem_2[428] <= 0;
    valid_1[429]  <=   0;valid_2[429]  <=   0;dirty_bit_1[429] <= 0;dirty_bit_2[429] <= 0;lru_counter_1[429] <= 0;lru_counter_2[429] <= 0;tag_1[429] <= 0;tag_2[429] <= 0;cache_mem_1[429] <= 0;cache_mem_2[429] <= 0;
    valid_1[430]  <=   0;valid_2[430]  <=   0;dirty_bit_1[430] <= 0;dirty_bit_2[430] <= 0;lru_counter_1[430] <= 0;lru_counter_2[430] <= 0;tag_1[430] <= 0;tag_2[430] <= 0;cache_mem_1[430] <= 0;cache_mem_2[430] <= 0;
    valid_1[431]  <=   0;valid_2[431]  <=   0;dirty_bit_1[431] <= 0;dirty_bit_2[431] <= 0;lru_counter_1[431] <= 0;lru_counter_2[431] <= 0;tag_1[431] <= 0;tag_2[431] <= 0;cache_mem_1[431] <= 0;cache_mem_2[431] <= 0;
    valid_1[432]  <=   0;valid_2[432]  <=   0;dirty_bit_1[432] <= 0;dirty_bit_2[432] <= 0;lru_counter_1[432] <= 0;lru_counter_2[432] <= 0;tag_1[432] <= 0;tag_2[432] <= 0;cache_mem_1[432] <= 0;cache_mem_2[432] <= 0;
    valid_1[433]  <=   0;valid_2[433]  <=   0;dirty_bit_1[433] <= 0;dirty_bit_2[433] <= 0;lru_counter_1[433] <= 0;lru_counter_2[433] <= 0;tag_1[433] <= 0;tag_2[433] <= 0;cache_mem_1[433] <= 0;cache_mem_2[433] <= 0;
    valid_1[434]  <=   0;valid_2[434]  <=   0;dirty_bit_1[434] <= 0;dirty_bit_2[434] <= 0;lru_counter_1[434] <= 0;lru_counter_2[434] <= 0;tag_1[434] <= 0;tag_2[434] <= 0;cache_mem_1[434] <= 0;cache_mem_2[434] <= 0;
    valid_1[435]  <=   0;valid_2[435]  <=   0;dirty_bit_1[435] <= 0;dirty_bit_2[435] <= 0;lru_counter_1[435] <= 0;lru_counter_2[435] <= 0;tag_1[435] <= 0;tag_2[435] <= 0;cache_mem_1[435] <= 0;cache_mem_2[435] <= 0;
    valid_1[436]  <=   0;valid_2[436]  <=   0;dirty_bit_1[436] <= 0;dirty_bit_2[436] <= 0;lru_counter_1[436] <= 0;lru_counter_2[436] <= 0;tag_1[436] <= 0;tag_2[436] <= 0;cache_mem_1[436] <= 0;cache_mem_2[436] <= 0;
    valid_1[437]  <=   0;valid_2[437]  <=   0;dirty_bit_1[437] <= 0;dirty_bit_2[437] <= 0;lru_counter_1[437] <= 0;lru_counter_2[437] <= 0;tag_1[437] <= 0;tag_2[437] <= 0;cache_mem_1[437] <= 0;cache_mem_2[437] <= 0;
    valid_1[438]  <=   0;valid_2[438]  <=   0;dirty_bit_1[438] <= 0;dirty_bit_2[438] <= 0;lru_counter_1[438] <= 0;lru_counter_2[438] <= 0;tag_1[438] <= 0;tag_2[438] <= 0;cache_mem_1[438] <= 0;cache_mem_2[438] <= 0;
    valid_1[439]  <=   0;valid_2[439]  <=   0;dirty_bit_1[439] <= 0;dirty_bit_2[439] <= 0;lru_counter_1[439] <= 0;lru_counter_2[439] <= 0;tag_1[439] <= 0;tag_2[439] <= 0;cache_mem_1[439] <= 0;cache_mem_2[439] <= 0;
    valid_1[440]  <=   0;valid_2[440]  <=   0;dirty_bit_1[440] <= 0;dirty_bit_2[440] <= 0;lru_counter_1[440] <= 0;lru_counter_2[440] <= 0;tag_1[440] <= 0;tag_2[440] <= 0;cache_mem_1[440] <= 0;cache_mem_2[440] <= 0;
    valid_1[441]  <=   0;valid_2[441]  <=   0;dirty_bit_1[441] <= 0;dirty_bit_2[441] <= 0;lru_counter_1[441] <= 0;lru_counter_2[441] <= 0;tag_1[441] <= 0;tag_2[441] <= 0;cache_mem_1[441] <= 0;cache_mem_2[441] <= 0;
    valid_1[442]  <=   0;valid_2[442]  <=   0;dirty_bit_1[442] <= 0;dirty_bit_2[442] <= 0;lru_counter_1[442] <= 0;lru_counter_2[442] <= 0;tag_1[442] <= 0;tag_2[442] <= 0;cache_mem_1[442] <= 0;cache_mem_2[442] <= 0;
    valid_1[443]  <=   0;valid_2[443]  <=   0;dirty_bit_1[443] <= 0;dirty_bit_2[443] <= 0;lru_counter_1[443] <= 0;lru_counter_2[443] <= 0;tag_1[443] <= 0;tag_2[443] <= 0;cache_mem_1[443] <= 0;cache_mem_2[443] <= 0;
    valid_1[444]  <=   0;valid_2[444]  <=   0;dirty_bit_1[444] <= 0;dirty_bit_2[444] <= 0;lru_counter_1[444] <= 0;lru_counter_2[444] <= 0;tag_1[444] <= 0;tag_2[444] <= 0;cache_mem_1[444] <= 0;cache_mem_2[444] <= 0;
    valid_1[445]  <=   0;valid_2[445]  <=   0;dirty_bit_1[445] <= 0;dirty_bit_2[445] <= 0;lru_counter_1[445] <= 0;lru_counter_2[445] <= 0;tag_1[445] <= 0;tag_2[445] <= 0;cache_mem_1[445] <= 0;cache_mem_2[445] <= 0;
    valid_1[446]  <=   0;valid_2[446]  <=   0;dirty_bit_1[446] <= 0;dirty_bit_2[446] <= 0;lru_counter_1[446] <= 0;lru_counter_2[446] <= 0;tag_1[446] <= 0;tag_2[446] <= 0;cache_mem_1[446] <= 0;cache_mem_2[446] <= 0;
    valid_1[447]  <=   0;valid_2[447]  <=   0;dirty_bit_1[447] <= 0;dirty_bit_2[447] <= 0;lru_counter_1[447] <= 0;lru_counter_2[447] <= 0;tag_1[447] <= 0;tag_2[447] <= 0;cache_mem_1[447] <= 0;cache_mem_2[447] <= 0;
    valid_1[448]  <=   0;valid_2[448]  <=   0;dirty_bit_1[448] <= 0;dirty_bit_2[448] <= 0;lru_counter_1[448] <= 0;lru_counter_2[448] <= 0;tag_1[448] <= 0;tag_2[448] <= 0;cache_mem_1[448] <= 0;cache_mem_2[448] <= 0;
    valid_1[449]  <=   0;valid_2[449]  <=   0;dirty_bit_1[449] <= 0;dirty_bit_2[449] <= 0;lru_counter_1[449] <= 0;lru_counter_2[449] <= 0;tag_1[449] <= 0;tag_2[449] <= 0;cache_mem_1[449] <= 0;cache_mem_2[449] <= 0;
    valid_1[450]  <=   0;valid_2[450]  <=   0;dirty_bit_1[450] <= 0;dirty_bit_2[450] <= 0;lru_counter_1[450] <= 0;lru_counter_2[450] <= 0;tag_1[450] <= 0;tag_2[450] <= 0;cache_mem_1[450] <= 0;cache_mem_2[450] <= 0;
    valid_1[451]  <=   0;valid_2[451]  <=   0;dirty_bit_1[451] <= 0;dirty_bit_2[451] <= 0;lru_counter_1[451] <= 0;lru_counter_2[451] <= 0;tag_1[451] <= 0;tag_2[451] <= 0;cache_mem_1[451] <= 0;cache_mem_2[451] <= 0;
    valid_1[452]  <=   0;valid_2[452]  <=   0;dirty_bit_1[452] <= 0;dirty_bit_2[452] <= 0;lru_counter_1[452] <= 0;lru_counter_2[452] <= 0;tag_1[452] <= 0;tag_2[452] <= 0;cache_mem_1[452] <= 0;cache_mem_2[452] <= 0;
    valid_1[453]  <=   0;valid_2[453]  <=   0;dirty_bit_1[453] <= 0;dirty_bit_2[453] <= 0;lru_counter_1[453] <= 0;lru_counter_2[453] <= 0;tag_1[453] <= 0;tag_2[453] <= 0;cache_mem_1[453] <= 0;cache_mem_2[453] <= 0;
    valid_1[454]  <=   0;valid_2[454]  <=   0;dirty_bit_1[454] <= 0;dirty_bit_2[454] <= 0;lru_counter_1[454] <= 0;lru_counter_2[454] <= 0;tag_1[454] <= 0;tag_2[454] <= 0;cache_mem_1[454] <= 0;cache_mem_2[454] <= 0;
    valid_1[455]  <=   0;valid_2[455]  <=   0;dirty_bit_1[455] <= 0;dirty_bit_2[455] <= 0;lru_counter_1[455] <= 0;lru_counter_2[455] <= 0;tag_1[455] <= 0;tag_2[455] <= 0;cache_mem_1[455] <= 0;cache_mem_2[455] <= 0;
    valid_1[456]  <=   0;valid_2[456]  <=   0;dirty_bit_1[456] <= 0;dirty_bit_2[456] <= 0;lru_counter_1[456] <= 0;lru_counter_2[456] <= 0;tag_1[456] <= 0;tag_2[456] <= 0;cache_mem_1[456] <= 0;cache_mem_2[456] <= 0;
    valid_1[457]  <=   0;valid_2[457]  <=   0;dirty_bit_1[457] <= 0;dirty_bit_2[457] <= 0;lru_counter_1[457] <= 0;lru_counter_2[457] <= 0;tag_1[457] <= 0;tag_2[457] <= 0;cache_mem_1[457] <= 0;cache_mem_2[457] <= 0;
    valid_1[458]  <=   0;valid_2[458]  <=   0;dirty_bit_1[458] <= 0;dirty_bit_2[458] <= 0;lru_counter_1[458] <= 0;lru_counter_2[458] <= 0;tag_1[458] <= 0;tag_2[458] <= 0;cache_mem_1[458] <= 0;cache_mem_2[458] <= 0;
    valid_1[459]  <=   0;valid_2[459]  <=   0;dirty_bit_1[459] <= 0;dirty_bit_2[459] <= 0;lru_counter_1[459] <= 0;lru_counter_2[459] <= 0;tag_1[459] <= 0;tag_2[459] <= 0;cache_mem_1[459] <= 0;cache_mem_2[459] <= 0;
    valid_1[460]  <=   0;valid_2[460]  <=   0;dirty_bit_1[460] <= 0;dirty_bit_2[460] <= 0;lru_counter_1[460] <= 0;lru_counter_2[460] <= 0;tag_1[460] <= 0;tag_2[460] <= 0;cache_mem_1[460] <= 0;cache_mem_2[460] <= 0;
    valid_1[461]  <=   0;valid_2[461]  <=   0;dirty_bit_1[461] <= 0;dirty_bit_2[461] <= 0;lru_counter_1[461] <= 0;lru_counter_2[461] <= 0;tag_1[461] <= 0;tag_2[461] <= 0;cache_mem_1[461] <= 0;cache_mem_2[461] <= 0;
    valid_1[462]  <=   0;valid_2[462]  <=   0;dirty_bit_1[462] <= 0;dirty_bit_2[462] <= 0;lru_counter_1[462] <= 0;lru_counter_2[462] <= 0;tag_1[462] <= 0;tag_2[462] <= 0;cache_mem_1[462] <= 0;cache_mem_2[462] <= 0;
    valid_1[463]  <=   0;valid_2[463]  <=   0;dirty_bit_1[463] <= 0;dirty_bit_2[463] <= 0;lru_counter_1[463] <= 0;lru_counter_2[463] <= 0;tag_1[463] <= 0;tag_2[463] <= 0;cache_mem_1[463] <= 0;cache_mem_2[463] <= 0;
    valid_1[464]  <=   0;valid_2[464]  <=   0;dirty_bit_1[464] <= 0;dirty_bit_2[464] <= 0;lru_counter_1[464] <= 0;lru_counter_2[464] <= 0;tag_1[464] <= 0;tag_2[464] <= 0;cache_mem_1[464] <= 0;cache_mem_2[464] <= 0;
    valid_1[465]  <=   0;valid_2[465]  <=   0;dirty_bit_1[465] <= 0;dirty_bit_2[465] <= 0;lru_counter_1[465] <= 0;lru_counter_2[465] <= 0;tag_1[465] <= 0;tag_2[465] <= 0;cache_mem_1[465] <= 0;cache_mem_2[465] <= 0;
    valid_1[466]  <=   0;valid_2[466]  <=   0;dirty_bit_1[466] <= 0;dirty_bit_2[466] <= 0;lru_counter_1[466] <= 0;lru_counter_2[466] <= 0;tag_1[466] <= 0;tag_2[466] <= 0;cache_mem_1[466] <= 0;cache_mem_2[466] <= 0;
    valid_1[467]  <=   0;valid_2[467]  <=   0;dirty_bit_1[467] <= 0;dirty_bit_2[467] <= 0;lru_counter_1[467] <= 0;lru_counter_2[467] <= 0;tag_1[467] <= 0;tag_2[467] <= 0;cache_mem_1[467] <= 0;cache_mem_2[467] <= 0;
    valid_1[468]  <=   0;valid_2[468]  <=   0;dirty_bit_1[468] <= 0;dirty_bit_2[468] <= 0;lru_counter_1[468] <= 0;lru_counter_2[468] <= 0;tag_1[468] <= 0;tag_2[468] <= 0;cache_mem_1[468] <= 0;cache_mem_2[468] <= 0;
    valid_1[469]  <=   0;valid_2[469]  <=   0;dirty_bit_1[469] <= 0;dirty_bit_2[469] <= 0;lru_counter_1[469] <= 0;lru_counter_2[469] <= 0;tag_1[469] <= 0;tag_2[469] <= 0;cache_mem_1[469] <= 0;cache_mem_2[469] <= 0;
    valid_1[470]  <=   0;valid_2[470]  <=   0;dirty_bit_1[470] <= 0;dirty_bit_2[470] <= 0;lru_counter_1[470] <= 0;lru_counter_2[470] <= 0;tag_1[470] <= 0;tag_2[470] <= 0;cache_mem_1[470] <= 0;cache_mem_2[470] <= 0;
    valid_1[471]  <=   0;valid_2[471]  <=   0;dirty_bit_1[471] <= 0;dirty_bit_2[471] <= 0;lru_counter_1[471] <= 0;lru_counter_2[471] <= 0;tag_1[471] <= 0;tag_2[471] <= 0;cache_mem_1[471] <= 0;cache_mem_2[471] <= 0;
    valid_1[472]  <=   0;valid_2[472]  <=   0;dirty_bit_1[472] <= 0;dirty_bit_2[472] <= 0;lru_counter_1[472] <= 0;lru_counter_2[472] <= 0;tag_1[472] <= 0;tag_2[472] <= 0;cache_mem_1[472] <= 0;cache_mem_2[472] <= 0;
    valid_1[473]  <=   0;valid_2[473]  <=   0;dirty_bit_1[473] <= 0;dirty_bit_2[473] <= 0;lru_counter_1[473] <= 0;lru_counter_2[473] <= 0;tag_1[473] <= 0;tag_2[473] <= 0;cache_mem_1[473] <= 0;cache_mem_2[473] <= 0;
    valid_1[474]  <=   0;valid_2[474]  <=   0;dirty_bit_1[474] <= 0;dirty_bit_2[474] <= 0;lru_counter_1[474] <= 0;lru_counter_2[474] <= 0;tag_1[474] <= 0;tag_2[474] <= 0;cache_mem_1[474] <= 0;cache_mem_2[474] <= 0;
    valid_1[475]  <=   0;valid_2[475]  <=   0;dirty_bit_1[475] <= 0;dirty_bit_2[475] <= 0;lru_counter_1[475] <= 0;lru_counter_2[475] <= 0;tag_1[475] <= 0;tag_2[475] <= 0;cache_mem_1[475] <= 0;cache_mem_2[475] <= 0;
    valid_1[476]  <=   0;valid_2[476]  <=   0;dirty_bit_1[476] <= 0;dirty_bit_2[476] <= 0;lru_counter_1[476] <= 0;lru_counter_2[476] <= 0;tag_1[476] <= 0;tag_2[476] <= 0;cache_mem_1[476] <= 0;cache_mem_2[476] <= 0;
    valid_1[477]  <=   0;valid_2[477]  <=   0;dirty_bit_1[477] <= 0;dirty_bit_2[477] <= 0;lru_counter_1[477] <= 0;lru_counter_2[477] <= 0;tag_1[477] <= 0;tag_2[477] <= 0;cache_mem_1[477] <= 0;cache_mem_2[477] <= 0;
    valid_1[478]  <=   0;valid_2[478]  <=   0;dirty_bit_1[478] <= 0;dirty_bit_2[478] <= 0;lru_counter_1[478] <= 0;lru_counter_2[478] <= 0;tag_1[478] <= 0;tag_2[478] <= 0;cache_mem_1[478] <= 0;cache_mem_2[478] <= 0;
    valid_1[479]  <=   0;valid_2[479]  <=   0;dirty_bit_1[479] <= 0;dirty_bit_2[479] <= 0;lru_counter_1[479] <= 0;lru_counter_2[479] <= 0;tag_1[479] <= 0;tag_2[479] <= 0;cache_mem_1[479] <= 0;cache_mem_2[479] <= 0;
    valid_1[480]  <=   0;valid_2[480]  <=   0;dirty_bit_1[480] <= 0;dirty_bit_2[480] <= 0;lru_counter_1[480] <= 0;lru_counter_2[480] <= 0;tag_1[480] <= 0;tag_2[480] <= 0;cache_mem_1[480] <= 0;cache_mem_2[480] <= 0;
    valid_1[481]  <=   0;valid_2[481]  <=   0;dirty_bit_1[481] <= 0;dirty_bit_2[481] <= 0;lru_counter_1[481] <= 0;lru_counter_2[481] <= 0;tag_1[481] <= 0;tag_2[481] <= 0;cache_mem_1[481] <= 0;cache_mem_2[481] <= 0;
    valid_1[482]  <=   0;valid_2[482]  <=   0;dirty_bit_1[482] <= 0;dirty_bit_2[482] <= 0;lru_counter_1[482] <= 0;lru_counter_2[482] <= 0;tag_1[482] <= 0;tag_2[482] <= 0;cache_mem_1[482] <= 0;cache_mem_2[482] <= 0;
    valid_1[483]  <=   0;valid_2[483]  <=   0;dirty_bit_1[483] <= 0;dirty_bit_2[483] <= 0;lru_counter_1[483] <= 0;lru_counter_2[483] <= 0;tag_1[483] <= 0;tag_2[483] <= 0;cache_mem_1[483] <= 0;cache_mem_2[483] <= 0;
    valid_1[484]  <=   0;valid_2[484]  <=   0;dirty_bit_1[484] <= 0;dirty_bit_2[484] <= 0;lru_counter_1[484] <= 0;lru_counter_2[484] <= 0;tag_1[484] <= 0;tag_2[484] <= 0;cache_mem_1[484] <= 0;cache_mem_2[484] <= 0;
    valid_1[485]  <=   0;valid_2[485]  <=   0;dirty_bit_1[485] <= 0;dirty_bit_2[485] <= 0;lru_counter_1[485] <= 0;lru_counter_2[485] <= 0;tag_1[485] <= 0;tag_2[485] <= 0;cache_mem_1[485] <= 0;cache_mem_2[485] <= 0;
    valid_1[486]  <=   0;valid_2[486]  <=   0;dirty_bit_1[486] <= 0;dirty_bit_2[486] <= 0;lru_counter_1[486] <= 0;lru_counter_2[486] <= 0;tag_1[486] <= 0;tag_2[486] <= 0;cache_mem_1[486] <= 0;cache_mem_2[486] <= 0;
    valid_1[487]  <=   0;valid_2[487]  <=   0;dirty_bit_1[487] <= 0;dirty_bit_2[487] <= 0;lru_counter_1[487] <= 0;lru_counter_2[487] <= 0;tag_1[487] <= 0;tag_2[487] <= 0;cache_mem_1[487] <= 0;cache_mem_2[487] <= 0;
    valid_1[488]  <=   0;valid_2[488]  <=   0;dirty_bit_1[488] <= 0;dirty_bit_2[488] <= 0;lru_counter_1[488] <= 0;lru_counter_2[488] <= 0;tag_1[488] <= 0;tag_2[488] <= 0;cache_mem_1[488] <= 0;cache_mem_2[488] <= 0;
    valid_1[489]  <=   0;valid_2[489]  <=   0;dirty_bit_1[489] <= 0;dirty_bit_2[489] <= 0;lru_counter_1[489] <= 0;lru_counter_2[489] <= 0;tag_1[489] <= 0;tag_2[489] <= 0;cache_mem_1[489] <= 0;cache_mem_2[489] <= 0;
    valid_1[490]  <=   0;valid_2[490]  <=   0;dirty_bit_1[490] <= 0;dirty_bit_2[490] <= 0;lru_counter_1[490] <= 0;lru_counter_2[490] <= 0;tag_1[490] <= 0;tag_2[490] <= 0;cache_mem_1[490] <= 0;cache_mem_2[490] <= 0;
    valid_1[491]  <=   0;valid_2[491]  <=   0;dirty_bit_1[491] <= 0;dirty_bit_2[491] <= 0;lru_counter_1[491] <= 0;lru_counter_2[491] <= 0;tag_1[491] <= 0;tag_2[491] <= 0;cache_mem_1[491] <= 0;cache_mem_2[491] <= 0;
    valid_1[492]  <=   0;valid_2[492]  <=   0;dirty_bit_1[492] <= 0;dirty_bit_2[492] <= 0;lru_counter_1[492] <= 0;lru_counter_2[492] <= 0;tag_1[492] <= 0;tag_2[492] <= 0;cache_mem_1[492] <= 0;cache_mem_2[492] <= 0;
    valid_1[493]  <=   0;valid_2[493]  <=   0;dirty_bit_1[493] <= 0;dirty_bit_2[493] <= 0;lru_counter_1[493] <= 0;lru_counter_2[493] <= 0;tag_1[493] <= 0;tag_2[493] <= 0;cache_mem_1[493] <= 0;cache_mem_2[493] <= 0;
    valid_1[494]  <=   0;valid_2[494]  <=   0;dirty_bit_1[494] <= 0;dirty_bit_2[494] <= 0;lru_counter_1[494] <= 0;lru_counter_2[494] <= 0;tag_1[494] <= 0;tag_2[494] <= 0;cache_mem_1[494] <= 0;cache_mem_2[494] <= 0;
    valid_1[495]  <=   0;valid_2[495]  <=   0;dirty_bit_1[495] <= 0;dirty_bit_2[495] <= 0;lru_counter_1[495] <= 0;lru_counter_2[495] <= 0;tag_1[495] <= 0;tag_2[495] <= 0;cache_mem_1[495] <= 0;cache_mem_2[495] <= 0;
    valid_1[496]  <=   0;valid_2[496]  <=   0;dirty_bit_1[496] <= 0;dirty_bit_2[496] <= 0;lru_counter_1[496] <= 0;lru_counter_2[496] <= 0;tag_1[496] <= 0;tag_2[496] <= 0;cache_mem_1[496] <= 0;cache_mem_2[496] <= 0;
    valid_1[497]  <=   0;valid_2[497]  <=   0;dirty_bit_1[497] <= 0;dirty_bit_2[497] <= 0;lru_counter_1[497] <= 0;lru_counter_2[497] <= 0;tag_1[497] <= 0;tag_2[497] <= 0;cache_mem_1[497] <= 0;cache_mem_2[497] <= 0;
    valid_1[498]  <=   0;valid_2[498]  <=   0;dirty_bit_1[498] <= 0;dirty_bit_2[498] <= 0;lru_counter_1[498] <= 0;lru_counter_2[498] <= 0;tag_1[498] <= 0;tag_2[498] <= 0;cache_mem_1[498] <= 0;cache_mem_2[498] <= 0;
    valid_1[499]  <=   0;valid_2[499]  <=   0;dirty_bit_1[499] <= 0;dirty_bit_2[499] <= 0;lru_counter_1[499] <= 0;lru_counter_2[499] <= 0;tag_1[499] <= 0;tag_2[499] <= 0;cache_mem_1[499] <= 0;cache_mem_2[499] <= 0;
    valid_1[500]  <=   0;valid_2[500]  <=   0;dirty_bit_1[500] <= 0;dirty_bit_2[500] <= 0;lru_counter_1[500] <= 0;lru_counter_2[500] <= 0;tag_1[500] <= 0;tag_2[500] <= 0;cache_mem_1[500] <= 0;cache_mem_2[500] <= 0;
    valid_1[501]  <=   0;valid_2[501]  <=   0;dirty_bit_1[501] <= 0;dirty_bit_2[501] <= 0;lru_counter_1[501] <= 0;lru_counter_2[501] <= 0;tag_1[501] <= 0;tag_2[501] <= 0;cache_mem_1[501] <= 0;cache_mem_2[501] <= 0;
    valid_1[502]  <=   0;valid_2[502]  <=   0;dirty_bit_1[502] <= 0;dirty_bit_2[502] <= 0;lru_counter_1[502] <= 0;lru_counter_2[502] <= 0;tag_1[502] <= 0;tag_2[502] <= 0;cache_mem_1[502] <= 0;cache_mem_2[502] <= 0;
    valid_1[503]  <=   0;valid_2[503]  <=   0;dirty_bit_1[503] <= 0;dirty_bit_2[503] <= 0;lru_counter_1[503] <= 0;lru_counter_2[503] <= 0;tag_1[503] <= 0;tag_2[503] <= 0;cache_mem_1[503] <= 0;cache_mem_2[503] <= 0;
    valid_1[504]  <=   0;valid_2[504]  <=   0;dirty_bit_1[504] <= 0;dirty_bit_2[504] <= 0;lru_counter_1[504] <= 0;lru_counter_2[504] <= 0;tag_1[504] <= 0;tag_2[504] <= 0;cache_mem_1[504] <= 0;cache_mem_2[504] <= 0;
    valid_1[505]  <=   0;valid_2[505]  <=   0;dirty_bit_1[505] <= 0;dirty_bit_2[505] <= 0;lru_counter_1[505] <= 0;lru_counter_2[505] <= 0;tag_1[505] <= 0;tag_2[505] <= 0;cache_mem_1[505] <= 0;cache_mem_2[505] <= 0;
    valid_1[506]  <=   0;valid_2[506]  <=   0;dirty_bit_1[506] <= 0;dirty_bit_2[506] <= 0;lru_counter_1[506] <= 0;lru_counter_2[506] <= 0;tag_1[506] <= 0;tag_2[506] <= 0;cache_mem_1[506] <= 0;cache_mem_2[506] <= 0;
    valid_1[507]  <=   0;valid_2[507]  <=   0;dirty_bit_1[507] <= 0;dirty_bit_2[507] <= 0;lru_counter_1[507] <= 0;lru_counter_2[507] <= 0;tag_1[507] <= 0;tag_2[507] <= 0;cache_mem_1[507] <= 0;cache_mem_2[507] <= 0;
    valid_1[508]  <=   0;valid_2[508]  <=   0;dirty_bit_1[508] <= 0;dirty_bit_2[508] <= 0;lru_counter_1[508] <= 0;lru_counter_2[508] <= 0;tag_1[508] <= 0;tag_2[508] <= 0;cache_mem_1[508] <= 0;cache_mem_2[508] <= 0;
    valid_1[509]  <=   0;valid_2[509]  <=   0;dirty_bit_1[509] <= 0;dirty_bit_2[509] <= 0;lru_counter_1[509] <= 0;lru_counter_2[509] <= 0;tag_1[509] <= 0;tag_2[509] <= 0;cache_mem_1[509] <= 0;cache_mem_2[509] <= 0;
    valid_1[510]  <=   0;valid_2[510]  <=   0;dirty_bit_1[510] <= 0;dirty_bit_2[510] <= 0;lru_counter_1[510] <= 0;lru_counter_2[510] <= 0;tag_1[510] <= 0;tag_2[510] <= 0;cache_mem_1[510] <= 0;cache_mem_2[510] <= 0;
    valid_1[511]  <=   0;valid_2[511]  <=   0;dirty_bit_1[511] <= 0;dirty_bit_2[511] <= 0;lru_counter_1[511] <= 0;lru_counter_2[511] <= 0;tag_1[511] <= 0;tag_2[511] <= 0;cache_mem_1[511] <= 0;cache_mem_2[511] <= 0;
    valid_1[512]  <=   0;valid_2[512]  <=   0;dirty_bit_1[512] <= 0;dirty_bit_2[512] <= 0;lru_counter_1[512] <= 0;lru_counter_2[512] <= 0;tag_1[512] <= 0;tag_2[512] <= 0;cache_mem_1[512] <= 0;cache_mem_2[512] <= 0;
    valid_1[513]  <=   0;valid_2[513]  <=   0;dirty_bit_1[513] <= 0;dirty_bit_2[513] <= 0;lru_counter_1[513] <= 0;lru_counter_2[513] <= 0;tag_1[513] <= 0;tag_2[513] <= 0;cache_mem_1[513] <= 0;cache_mem_2[513] <= 0;
    valid_1[514]  <=   0;valid_2[514]  <=   0;dirty_bit_1[514] <= 0;dirty_bit_2[514] <= 0;lru_counter_1[514] <= 0;lru_counter_2[514] <= 0;tag_1[514] <= 0;tag_2[514] <= 0;cache_mem_1[514] <= 0;cache_mem_2[514] <= 0;
    valid_1[515]  <=   0;valid_2[515]  <=   0;dirty_bit_1[515] <= 0;dirty_bit_2[515] <= 0;lru_counter_1[515] <= 0;lru_counter_2[515] <= 0;tag_1[515] <= 0;tag_2[515] <= 0;cache_mem_1[515] <= 0;cache_mem_2[515] <= 0;
    valid_1[516]  <=   0;valid_2[516]  <=   0;dirty_bit_1[516] <= 0;dirty_bit_2[516] <= 0;lru_counter_1[516] <= 0;lru_counter_2[516] <= 0;tag_1[516] <= 0;tag_2[516] <= 0;cache_mem_1[516] <= 0;cache_mem_2[516] <= 0;
    valid_1[517]  <=   0;valid_2[517]  <=   0;dirty_bit_1[517] <= 0;dirty_bit_2[517] <= 0;lru_counter_1[517] <= 0;lru_counter_2[517] <= 0;tag_1[517] <= 0;tag_2[517] <= 0;cache_mem_1[517] <= 0;cache_mem_2[517] <= 0;
    valid_1[518]  <=   0;valid_2[518]  <=   0;dirty_bit_1[518] <= 0;dirty_bit_2[518] <= 0;lru_counter_1[518] <= 0;lru_counter_2[518] <= 0;tag_1[518] <= 0;tag_2[518] <= 0;cache_mem_1[518] <= 0;cache_mem_2[518] <= 0;
    valid_1[519]  <=   0;valid_2[519]  <=   0;dirty_bit_1[519] <= 0;dirty_bit_2[519] <= 0;lru_counter_1[519] <= 0;lru_counter_2[519] <= 0;tag_1[519] <= 0;tag_2[519] <= 0;cache_mem_1[519] <= 0;cache_mem_2[519] <= 0;
    valid_1[520]  <=   0;valid_2[520]  <=   0;dirty_bit_1[520] <= 0;dirty_bit_2[520] <= 0;lru_counter_1[520] <= 0;lru_counter_2[520] <= 0;tag_1[520] <= 0;tag_2[520] <= 0;cache_mem_1[520] <= 0;cache_mem_2[520] <= 0;
    valid_1[521]  <=   0;valid_2[521]  <=   0;dirty_bit_1[521] <= 0;dirty_bit_2[521] <= 0;lru_counter_1[521] <= 0;lru_counter_2[521] <= 0;tag_1[521] <= 0;tag_2[521] <= 0;cache_mem_1[521] <= 0;cache_mem_2[521] <= 0;
    valid_1[522]  <=   0;valid_2[522]  <=   0;dirty_bit_1[522] <= 0;dirty_bit_2[522] <= 0;lru_counter_1[522] <= 0;lru_counter_2[522] <= 0;tag_1[522] <= 0;tag_2[522] <= 0;cache_mem_1[522] <= 0;cache_mem_2[522] <= 0;
    valid_1[523]  <=   0;valid_2[523]  <=   0;dirty_bit_1[523] <= 0;dirty_bit_2[523] <= 0;lru_counter_1[523] <= 0;lru_counter_2[523] <= 0;tag_1[523] <= 0;tag_2[523] <= 0;cache_mem_1[523] <= 0;cache_mem_2[523] <= 0;
    valid_1[524]  <=   0;valid_2[524]  <=   0;dirty_bit_1[524] <= 0;dirty_bit_2[524] <= 0;lru_counter_1[524] <= 0;lru_counter_2[524] <= 0;tag_1[524] <= 0;tag_2[524] <= 0;cache_mem_1[524] <= 0;cache_mem_2[524] <= 0;
    valid_1[525]  <=   0;valid_2[525]  <=   0;dirty_bit_1[525] <= 0;dirty_bit_2[525] <= 0;lru_counter_1[525] <= 0;lru_counter_2[525] <= 0;tag_1[525] <= 0;tag_2[525] <= 0;cache_mem_1[525] <= 0;cache_mem_2[525] <= 0;
    valid_1[526]  <=   0;valid_2[526]  <=   0;dirty_bit_1[526] <= 0;dirty_bit_2[526] <= 0;lru_counter_1[526] <= 0;lru_counter_2[526] <= 0;tag_1[526] <= 0;tag_2[526] <= 0;cache_mem_1[526] <= 0;cache_mem_2[526] <= 0;
    valid_1[527]  <=   0;valid_2[527]  <=   0;dirty_bit_1[527] <= 0;dirty_bit_2[527] <= 0;lru_counter_1[527] <= 0;lru_counter_2[527] <= 0;tag_1[527] <= 0;tag_2[527] <= 0;cache_mem_1[527] <= 0;cache_mem_2[527] <= 0;
    valid_1[528]  <=   0;valid_2[528]  <=   0;dirty_bit_1[528] <= 0;dirty_bit_2[528] <= 0;lru_counter_1[528] <= 0;lru_counter_2[528] <= 0;tag_1[528] <= 0;tag_2[528] <= 0;cache_mem_1[528] <= 0;cache_mem_2[528] <= 0;
    valid_1[529]  <=   0;valid_2[529]  <=   0;dirty_bit_1[529] <= 0;dirty_bit_2[529] <= 0;lru_counter_1[529] <= 0;lru_counter_2[529] <= 0;tag_1[529] <= 0;tag_2[529] <= 0;cache_mem_1[529] <= 0;cache_mem_2[529] <= 0;
    valid_1[530]  <=   0;valid_2[530]  <=   0;dirty_bit_1[530] <= 0;dirty_bit_2[530] <= 0;lru_counter_1[530] <= 0;lru_counter_2[530] <= 0;tag_1[530] <= 0;tag_2[530] <= 0;cache_mem_1[530] <= 0;cache_mem_2[530] <= 0;
    valid_1[531]  <=   0;valid_2[531]  <=   0;dirty_bit_1[531] <= 0;dirty_bit_2[531] <= 0;lru_counter_1[531] <= 0;lru_counter_2[531] <= 0;tag_1[531] <= 0;tag_2[531] <= 0;cache_mem_1[531] <= 0;cache_mem_2[531] <= 0;
    valid_1[532]  <=   0;valid_2[532]  <=   0;dirty_bit_1[532] <= 0;dirty_bit_2[532] <= 0;lru_counter_1[532] <= 0;lru_counter_2[532] <= 0;tag_1[532] <= 0;tag_2[532] <= 0;cache_mem_1[532] <= 0;cache_mem_2[532] <= 0;
    valid_1[533]  <=   0;valid_2[533]  <=   0;dirty_bit_1[533] <= 0;dirty_bit_2[533] <= 0;lru_counter_1[533] <= 0;lru_counter_2[533] <= 0;tag_1[533] <= 0;tag_2[533] <= 0;cache_mem_1[533] <= 0;cache_mem_2[533] <= 0;
    valid_1[534]  <=   0;valid_2[534]  <=   0;dirty_bit_1[534] <= 0;dirty_bit_2[534] <= 0;lru_counter_1[534] <= 0;lru_counter_2[534] <= 0;tag_1[534] <= 0;tag_2[534] <= 0;cache_mem_1[534] <= 0;cache_mem_2[534] <= 0;
    valid_1[535]  <=   0;valid_2[535]  <=   0;dirty_bit_1[535] <= 0;dirty_bit_2[535] <= 0;lru_counter_1[535] <= 0;lru_counter_2[535] <= 0;tag_1[535] <= 0;tag_2[535] <= 0;cache_mem_1[535] <= 0;cache_mem_2[535] <= 0;
    valid_1[536]  <=   0;valid_2[536]  <=   0;dirty_bit_1[536] <= 0;dirty_bit_2[536] <= 0;lru_counter_1[536] <= 0;lru_counter_2[536] <= 0;tag_1[536] <= 0;tag_2[536] <= 0;cache_mem_1[536] <= 0;cache_mem_2[536] <= 0;
    valid_1[537]  <=   0;valid_2[537]  <=   0;dirty_bit_1[537] <= 0;dirty_bit_2[537] <= 0;lru_counter_1[537] <= 0;lru_counter_2[537] <= 0;tag_1[537] <= 0;tag_2[537] <= 0;cache_mem_1[537] <= 0;cache_mem_2[537] <= 0;
    valid_1[538]  <=   0;valid_2[538]  <=   0;dirty_bit_1[538] <= 0;dirty_bit_2[538] <= 0;lru_counter_1[538] <= 0;lru_counter_2[538] <= 0;tag_1[538] <= 0;tag_2[538] <= 0;cache_mem_1[538] <= 0;cache_mem_2[538] <= 0;
    valid_1[539]  <=   0;valid_2[539]  <=   0;dirty_bit_1[539] <= 0;dirty_bit_2[539] <= 0;lru_counter_1[539] <= 0;lru_counter_2[539] <= 0;tag_1[539] <= 0;tag_2[539] <= 0;cache_mem_1[539] <= 0;cache_mem_2[539] <= 0;
    valid_1[540]  <=   0;valid_2[540]  <=   0;dirty_bit_1[540] <= 0;dirty_bit_2[540] <= 0;lru_counter_1[540] <= 0;lru_counter_2[540] <= 0;tag_1[540] <= 0;tag_2[540] <= 0;cache_mem_1[540] <= 0;cache_mem_2[540] <= 0;
    valid_1[541]  <=   0;valid_2[541]  <=   0;dirty_bit_1[541] <= 0;dirty_bit_2[541] <= 0;lru_counter_1[541] <= 0;lru_counter_2[541] <= 0;tag_1[541] <= 0;tag_2[541] <= 0;cache_mem_1[541] <= 0;cache_mem_2[541] <= 0;
    valid_1[542]  <=   0;valid_2[542]  <=   0;dirty_bit_1[542] <= 0;dirty_bit_2[542] <= 0;lru_counter_1[542] <= 0;lru_counter_2[542] <= 0;tag_1[542] <= 0;tag_2[542] <= 0;cache_mem_1[542] <= 0;cache_mem_2[542] <= 0;
    valid_1[543]  <=   0;valid_2[543]  <=   0;dirty_bit_1[543] <= 0;dirty_bit_2[543] <= 0;lru_counter_1[543] <= 0;lru_counter_2[543] <= 0;tag_1[543] <= 0;tag_2[543] <= 0;cache_mem_1[543] <= 0;cache_mem_2[543] <= 0;
    valid_1[544]  <=   0;valid_2[544]  <=   0;dirty_bit_1[544] <= 0;dirty_bit_2[544] <= 0;lru_counter_1[544] <= 0;lru_counter_2[544] <= 0;tag_1[544] <= 0;tag_2[544] <= 0;cache_mem_1[544] <= 0;cache_mem_2[544] <= 0;
    valid_1[545]  <=   0;valid_2[545]  <=   0;dirty_bit_1[545] <= 0;dirty_bit_2[545] <= 0;lru_counter_1[545] <= 0;lru_counter_2[545] <= 0;tag_1[545] <= 0;tag_2[545] <= 0;cache_mem_1[545] <= 0;cache_mem_2[545] <= 0;
    valid_1[546]  <=   0;valid_2[546]  <=   0;dirty_bit_1[546] <= 0;dirty_bit_2[546] <= 0;lru_counter_1[546] <= 0;lru_counter_2[546] <= 0;tag_1[546] <= 0;tag_2[546] <= 0;cache_mem_1[546] <= 0;cache_mem_2[546] <= 0;
    valid_1[547]  <=   0;valid_2[547]  <=   0;dirty_bit_1[547] <= 0;dirty_bit_2[547] <= 0;lru_counter_1[547] <= 0;lru_counter_2[547] <= 0;tag_1[547] <= 0;tag_2[547] <= 0;cache_mem_1[547] <= 0;cache_mem_2[547] <= 0;
    valid_1[548]  <=   0;valid_2[548]  <=   0;dirty_bit_1[548] <= 0;dirty_bit_2[548] <= 0;lru_counter_1[548] <= 0;lru_counter_2[548] <= 0;tag_1[548] <= 0;tag_2[548] <= 0;cache_mem_1[548] <= 0;cache_mem_2[548] <= 0;
    valid_1[549]  <=   0;valid_2[549]  <=   0;dirty_bit_1[549] <= 0;dirty_bit_2[549] <= 0;lru_counter_1[549] <= 0;lru_counter_2[549] <= 0;tag_1[549] <= 0;tag_2[549] <= 0;cache_mem_1[549] <= 0;cache_mem_2[549] <= 0;
    valid_1[550]  <=   0;valid_2[550]  <=   0;dirty_bit_1[550] <= 0;dirty_bit_2[550] <= 0;lru_counter_1[550] <= 0;lru_counter_2[550] <= 0;tag_1[550] <= 0;tag_2[550] <= 0;cache_mem_1[550] <= 0;cache_mem_2[550] <= 0;
    valid_1[551]  <=   0;valid_2[551]  <=   0;dirty_bit_1[551] <= 0;dirty_bit_2[551] <= 0;lru_counter_1[551] <= 0;lru_counter_2[551] <= 0;tag_1[551] <= 0;tag_2[551] <= 0;cache_mem_1[551] <= 0;cache_mem_2[551] <= 0;
    valid_1[552]  <=   0;valid_2[552]  <=   0;dirty_bit_1[552] <= 0;dirty_bit_2[552] <= 0;lru_counter_1[552] <= 0;lru_counter_2[552] <= 0;tag_1[552] <= 0;tag_2[552] <= 0;cache_mem_1[552] <= 0;cache_mem_2[552] <= 0;
    valid_1[553]  <=   0;valid_2[553]  <=   0;dirty_bit_1[553] <= 0;dirty_bit_2[553] <= 0;lru_counter_1[553] <= 0;lru_counter_2[553] <= 0;tag_1[553] <= 0;tag_2[553] <= 0;cache_mem_1[553] <= 0;cache_mem_2[553] <= 0;
    valid_1[554]  <=   0;valid_2[554]  <=   0;dirty_bit_1[554] <= 0;dirty_bit_2[554] <= 0;lru_counter_1[554] <= 0;lru_counter_2[554] <= 0;tag_1[554] <= 0;tag_2[554] <= 0;cache_mem_1[554] <= 0;cache_mem_2[554] <= 0;
    valid_1[555]  <=   0;valid_2[555]  <=   0;dirty_bit_1[555] <= 0;dirty_bit_2[555] <= 0;lru_counter_1[555] <= 0;lru_counter_2[555] <= 0;tag_1[555] <= 0;tag_2[555] <= 0;cache_mem_1[555] <= 0;cache_mem_2[555] <= 0;
    valid_1[556]  <=   0;valid_2[556]  <=   0;dirty_bit_1[556] <= 0;dirty_bit_2[556] <= 0;lru_counter_1[556] <= 0;lru_counter_2[556] <= 0;tag_1[556] <= 0;tag_2[556] <= 0;cache_mem_1[556] <= 0;cache_mem_2[556] <= 0;
    valid_1[557]  <=   0;valid_2[557]  <=   0;dirty_bit_1[557] <= 0;dirty_bit_2[557] <= 0;lru_counter_1[557] <= 0;lru_counter_2[557] <= 0;tag_1[557] <= 0;tag_2[557] <= 0;cache_mem_1[557] <= 0;cache_mem_2[557] <= 0;
    valid_1[558]  <=   0;valid_2[558]  <=   0;dirty_bit_1[558] <= 0;dirty_bit_2[558] <= 0;lru_counter_1[558] <= 0;lru_counter_2[558] <= 0;tag_1[558] <= 0;tag_2[558] <= 0;cache_mem_1[558] <= 0;cache_mem_2[558] <= 0;
    valid_1[559]  <=   0;valid_2[559]  <=   0;dirty_bit_1[559] <= 0;dirty_bit_2[559] <= 0;lru_counter_1[559] <= 0;lru_counter_2[559] <= 0;tag_1[559] <= 0;tag_2[559] <= 0;cache_mem_1[559] <= 0;cache_mem_2[559] <= 0;
    valid_1[560]  <=   0;valid_2[560]  <=   0;dirty_bit_1[560] <= 0;dirty_bit_2[560] <= 0;lru_counter_1[560] <= 0;lru_counter_2[560] <= 0;tag_1[560] <= 0;tag_2[560] <= 0;cache_mem_1[560] <= 0;cache_mem_2[560] <= 0;
    valid_1[561]  <=   0;valid_2[561]  <=   0;dirty_bit_1[561] <= 0;dirty_bit_2[561] <= 0;lru_counter_1[561] <= 0;lru_counter_2[561] <= 0;tag_1[561] <= 0;tag_2[561] <= 0;cache_mem_1[561] <= 0;cache_mem_2[561] <= 0;
    valid_1[562]  <=   0;valid_2[562]  <=   0;dirty_bit_1[562] <= 0;dirty_bit_2[562] <= 0;lru_counter_1[562] <= 0;lru_counter_2[562] <= 0;tag_1[562] <= 0;tag_2[562] <= 0;cache_mem_1[562] <= 0;cache_mem_2[562] <= 0;
    valid_1[563]  <=   0;valid_2[563]  <=   0;dirty_bit_1[563] <= 0;dirty_bit_2[563] <= 0;lru_counter_1[563] <= 0;lru_counter_2[563] <= 0;tag_1[563] <= 0;tag_2[563] <= 0;cache_mem_1[563] <= 0;cache_mem_2[563] <= 0;
    valid_1[564]  <=   0;valid_2[564]  <=   0;dirty_bit_1[564] <= 0;dirty_bit_2[564] <= 0;lru_counter_1[564] <= 0;lru_counter_2[564] <= 0;tag_1[564] <= 0;tag_2[564] <= 0;cache_mem_1[564] <= 0;cache_mem_2[564] <= 0;
    valid_1[565]  <=   0;valid_2[565]  <=   0;dirty_bit_1[565] <= 0;dirty_bit_2[565] <= 0;lru_counter_1[565] <= 0;lru_counter_2[565] <= 0;tag_1[565] <= 0;tag_2[565] <= 0;cache_mem_1[565] <= 0;cache_mem_2[565] <= 0;
    valid_1[566]  <=   0;valid_2[566]  <=   0;dirty_bit_1[566] <= 0;dirty_bit_2[566] <= 0;lru_counter_1[566] <= 0;lru_counter_2[566] <= 0;tag_1[566] <= 0;tag_2[566] <= 0;cache_mem_1[566] <= 0;cache_mem_2[566] <= 0;
    valid_1[567]  <=   0;valid_2[567]  <=   0;dirty_bit_1[567] <= 0;dirty_bit_2[567] <= 0;lru_counter_1[567] <= 0;lru_counter_2[567] <= 0;tag_1[567] <= 0;tag_2[567] <= 0;cache_mem_1[567] <= 0;cache_mem_2[567] <= 0;
    valid_1[568]  <=   0;valid_2[568]  <=   0;dirty_bit_1[568] <= 0;dirty_bit_2[568] <= 0;lru_counter_1[568] <= 0;lru_counter_2[568] <= 0;tag_1[568] <= 0;tag_2[568] <= 0;cache_mem_1[568] <= 0;cache_mem_2[568] <= 0;
    valid_1[569]  <=   0;valid_2[569]  <=   0;dirty_bit_1[569] <= 0;dirty_bit_2[569] <= 0;lru_counter_1[569] <= 0;lru_counter_2[569] <= 0;tag_1[569] <= 0;tag_2[569] <= 0;cache_mem_1[569] <= 0;cache_mem_2[569] <= 0;
    valid_1[570]  <=   0;valid_2[570]  <=   0;dirty_bit_1[570] <= 0;dirty_bit_2[570] <= 0;lru_counter_1[570] <= 0;lru_counter_2[570] <= 0;tag_1[570] <= 0;tag_2[570] <= 0;cache_mem_1[570] <= 0;cache_mem_2[570] <= 0;
    valid_1[571]  <=   0;valid_2[571]  <=   0;dirty_bit_1[571] <= 0;dirty_bit_2[571] <= 0;lru_counter_1[571] <= 0;lru_counter_2[571] <= 0;tag_1[571] <= 0;tag_2[571] <= 0;cache_mem_1[571] <= 0;cache_mem_2[571] <= 0;
    valid_1[572]  <=   0;valid_2[572]  <=   0;dirty_bit_1[572] <= 0;dirty_bit_2[572] <= 0;lru_counter_1[572] <= 0;lru_counter_2[572] <= 0;tag_1[572] <= 0;tag_2[572] <= 0;cache_mem_1[572] <= 0;cache_mem_2[572] <= 0;
    valid_1[573]  <=   0;valid_2[573]  <=   0;dirty_bit_1[573] <= 0;dirty_bit_2[573] <= 0;lru_counter_1[573] <= 0;lru_counter_2[573] <= 0;tag_1[573] <= 0;tag_2[573] <= 0;cache_mem_1[573] <= 0;cache_mem_2[573] <= 0;
    valid_1[574]  <=   0;valid_2[574]  <=   0;dirty_bit_1[574] <= 0;dirty_bit_2[574] <= 0;lru_counter_1[574] <= 0;lru_counter_2[574] <= 0;tag_1[574] <= 0;tag_2[574] <= 0;cache_mem_1[574] <= 0;cache_mem_2[574] <= 0;
    valid_1[575]  <=   0;valid_2[575]  <=   0;dirty_bit_1[575] <= 0;dirty_bit_2[575] <= 0;lru_counter_1[575] <= 0;lru_counter_2[575] <= 0;tag_1[575] <= 0;tag_2[575] <= 0;cache_mem_1[575] <= 0;cache_mem_2[575] <= 0;
    valid_1[576]  <=   0;valid_2[576]  <=   0;dirty_bit_1[576] <= 0;dirty_bit_2[576] <= 0;lru_counter_1[576] <= 0;lru_counter_2[576] <= 0;tag_1[576] <= 0;tag_2[576] <= 0;cache_mem_1[576] <= 0;cache_mem_2[576] <= 0;
    valid_1[577]  <=   0;valid_2[577]  <=   0;dirty_bit_1[577] <= 0;dirty_bit_2[577] <= 0;lru_counter_1[577] <= 0;lru_counter_2[577] <= 0;tag_1[577] <= 0;tag_2[577] <= 0;cache_mem_1[577] <= 0;cache_mem_2[577] <= 0;
    valid_1[578]  <=   0;valid_2[578]  <=   0;dirty_bit_1[578] <= 0;dirty_bit_2[578] <= 0;lru_counter_1[578] <= 0;lru_counter_2[578] <= 0;tag_1[578] <= 0;tag_2[578] <= 0;cache_mem_1[578] <= 0;cache_mem_2[578] <= 0;
    valid_1[579]  <=   0;valid_2[579]  <=   0;dirty_bit_1[579] <= 0;dirty_bit_2[579] <= 0;lru_counter_1[579] <= 0;lru_counter_2[579] <= 0;tag_1[579] <= 0;tag_2[579] <= 0;cache_mem_1[579] <= 0;cache_mem_2[579] <= 0;
    valid_1[580]  <=   0;valid_2[580]  <=   0;dirty_bit_1[580] <= 0;dirty_bit_2[580] <= 0;lru_counter_1[580] <= 0;lru_counter_2[580] <= 0;tag_1[580] <= 0;tag_2[580] <= 0;cache_mem_1[580] <= 0;cache_mem_2[580] <= 0;
    valid_1[581]  <=   0;valid_2[581]  <=   0;dirty_bit_1[581] <= 0;dirty_bit_2[581] <= 0;lru_counter_1[581] <= 0;lru_counter_2[581] <= 0;tag_1[581] <= 0;tag_2[581] <= 0;cache_mem_1[581] <= 0;cache_mem_2[581] <= 0;
    valid_1[582]  <=   0;valid_2[582]  <=   0;dirty_bit_1[582] <= 0;dirty_bit_2[582] <= 0;lru_counter_1[582] <= 0;lru_counter_2[582] <= 0;tag_1[582] <= 0;tag_2[582] <= 0;cache_mem_1[582] <= 0;cache_mem_2[582] <= 0;
    valid_1[583]  <=   0;valid_2[583]  <=   0;dirty_bit_1[583] <= 0;dirty_bit_2[583] <= 0;lru_counter_1[583] <= 0;lru_counter_2[583] <= 0;tag_1[583] <= 0;tag_2[583] <= 0;cache_mem_1[583] <= 0;cache_mem_2[583] <= 0;
    valid_1[584]  <=   0;valid_2[584]  <=   0;dirty_bit_1[584] <= 0;dirty_bit_2[584] <= 0;lru_counter_1[584] <= 0;lru_counter_2[584] <= 0;tag_1[584] <= 0;tag_2[584] <= 0;cache_mem_1[584] <= 0;cache_mem_2[584] <= 0;
    valid_1[585]  <=   0;valid_2[585]  <=   0;dirty_bit_1[585] <= 0;dirty_bit_2[585] <= 0;lru_counter_1[585] <= 0;lru_counter_2[585] <= 0;tag_1[585] <= 0;tag_2[585] <= 0;cache_mem_1[585] <= 0;cache_mem_2[585] <= 0;
    valid_1[586]  <=   0;valid_2[586]  <=   0;dirty_bit_1[586] <= 0;dirty_bit_2[586] <= 0;lru_counter_1[586] <= 0;lru_counter_2[586] <= 0;tag_1[586] <= 0;tag_2[586] <= 0;cache_mem_1[586] <= 0;cache_mem_2[586] <= 0;
    valid_1[587]  <=   0;valid_2[587]  <=   0;dirty_bit_1[587] <= 0;dirty_bit_2[587] <= 0;lru_counter_1[587] <= 0;lru_counter_2[587] <= 0;tag_1[587] <= 0;tag_2[587] <= 0;cache_mem_1[587] <= 0;cache_mem_2[587] <= 0;
    valid_1[588]  <=   0;valid_2[588]  <=   0;dirty_bit_1[588] <= 0;dirty_bit_2[588] <= 0;lru_counter_1[588] <= 0;lru_counter_2[588] <= 0;tag_1[588] <= 0;tag_2[588] <= 0;cache_mem_1[588] <= 0;cache_mem_2[588] <= 0;
    valid_1[589]  <=   0;valid_2[589]  <=   0;dirty_bit_1[589] <= 0;dirty_bit_2[589] <= 0;lru_counter_1[589] <= 0;lru_counter_2[589] <= 0;tag_1[589] <= 0;tag_2[589] <= 0;cache_mem_1[589] <= 0;cache_mem_2[589] <= 0;
    valid_1[590]  <=   0;valid_2[590]  <=   0;dirty_bit_1[590] <= 0;dirty_bit_2[590] <= 0;lru_counter_1[590] <= 0;lru_counter_2[590] <= 0;tag_1[590] <= 0;tag_2[590] <= 0;cache_mem_1[590] <= 0;cache_mem_2[590] <= 0;
    valid_1[591]  <=   0;valid_2[591]  <=   0;dirty_bit_1[591] <= 0;dirty_bit_2[591] <= 0;lru_counter_1[591] <= 0;lru_counter_2[591] <= 0;tag_1[591] <= 0;tag_2[591] <= 0;cache_mem_1[591] <= 0;cache_mem_2[591] <= 0;
    valid_1[592]  <=   0;valid_2[592]  <=   0;dirty_bit_1[592] <= 0;dirty_bit_2[592] <= 0;lru_counter_1[592] <= 0;lru_counter_2[592] <= 0;tag_1[592] <= 0;tag_2[592] <= 0;cache_mem_1[592] <= 0;cache_mem_2[592] <= 0;
    valid_1[593]  <=   0;valid_2[593]  <=   0;dirty_bit_1[593] <= 0;dirty_bit_2[593] <= 0;lru_counter_1[593] <= 0;lru_counter_2[593] <= 0;tag_1[593] <= 0;tag_2[593] <= 0;cache_mem_1[593] <= 0;cache_mem_2[593] <= 0;
    valid_1[594]  <=   0;valid_2[594]  <=   0;dirty_bit_1[594] <= 0;dirty_bit_2[594] <= 0;lru_counter_1[594] <= 0;lru_counter_2[594] <= 0;tag_1[594] <= 0;tag_2[594] <= 0;cache_mem_1[594] <= 0;cache_mem_2[594] <= 0;
    valid_1[595]  <=   0;valid_2[595]  <=   0;dirty_bit_1[595] <= 0;dirty_bit_2[595] <= 0;lru_counter_1[595] <= 0;lru_counter_2[595] <= 0;tag_1[595] <= 0;tag_2[595] <= 0;cache_mem_1[595] <= 0;cache_mem_2[595] <= 0;
    valid_1[596]  <=   0;valid_2[596]  <=   0;dirty_bit_1[596] <= 0;dirty_bit_2[596] <= 0;lru_counter_1[596] <= 0;lru_counter_2[596] <= 0;tag_1[596] <= 0;tag_2[596] <= 0;cache_mem_1[596] <= 0;cache_mem_2[596] <= 0;
    valid_1[597]  <=   0;valid_2[597]  <=   0;dirty_bit_1[597] <= 0;dirty_bit_2[597] <= 0;lru_counter_1[597] <= 0;lru_counter_2[597] <= 0;tag_1[597] <= 0;tag_2[597] <= 0;cache_mem_1[597] <= 0;cache_mem_2[597] <= 0;
    valid_1[598]  <=   0;valid_2[598]  <=   0;dirty_bit_1[598] <= 0;dirty_bit_2[598] <= 0;lru_counter_1[598] <= 0;lru_counter_2[598] <= 0;tag_1[598] <= 0;tag_2[598] <= 0;cache_mem_1[598] <= 0;cache_mem_2[598] <= 0;
    valid_1[599]  <=   0;valid_2[599]  <=   0;dirty_bit_1[599] <= 0;dirty_bit_2[599] <= 0;lru_counter_1[599] <= 0;lru_counter_2[599] <= 0;tag_1[599] <= 0;tag_2[599] <= 0;cache_mem_1[599] <= 0;cache_mem_2[599] <= 0;
    valid_1[600]  <=   0;valid_2[600]  <=   0;dirty_bit_1[600] <= 0;dirty_bit_2[600] <= 0;lru_counter_1[600] <= 0;lru_counter_2[600] <= 0;tag_1[600] <= 0;tag_2[600] <= 0;cache_mem_1[600] <= 0;cache_mem_2[600] <= 0;
    valid_1[601]  <=   0;valid_2[601]  <=   0;dirty_bit_1[601] <= 0;dirty_bit_2[601] <= 0;lru_counter_1[601] <= 0;lru_counter_2[601] <= 0;tag_1[601] <= 0;tag_2[601] <= 0;cache_mem_1[601] <= 0;cache_mem_2[601] <= 0;
    valid_1[602]  <=   0;valid_2[602]  <=   0;dirty_bit_1[602] <= 0;dirty_bit_2[602] <= 0;lru_counter_1[602] <= 0;lru_counter_2[602] <= 0;tag_1[602] <= 0;tag_2[602] <= 0;cache_mem_1[602] <= 0;cache_mem_2[602] <= 0;
    valid_1[603]  <=   0;valid_2[603]  <=   0;dirty_bit_1[603] <= 0;dirty_bit_2[603] <= 0;lru_counter_1[603] <= 0;lru_counter_2[603] <= 0;tag_1[603] <= 0;tag_2[603] <= 0;cache_mem_1[603] <= 0;cache_mem_2[603] <= 0;
    valid_1[604]  <=   0;valid_2[604]  <=   0;dirty_bit_1[604] <= 0;dirty_bit_2[604] <= 0;lru_counter_1[604] <= 0;lru_counter_2[604] <= 0;tag_1[604] <= 0;tag_2[604] <= 0;cache_mem_1[604] <= 0;cache_mem_2[604] <= 0;
    valid_1[605]  <=   0;valid_2[605]  <=   0;dirty_bit_1[605] <= 0;dirty_bit_2[605] <= 0;lru_counter_1[605] <= 0;lru_counter_2[605] <= 0;tag_1[605] <= 0;tag_2[605] <= 0;cache_mem_1[605] <= 0;cache_mem_2[605] <= 0;
    valid_1[606]  <=   0;valid_2[606]  <=   0;dirty_bit_1[606] <= 0;dirty_bit_2[606] <= 0;lru_counter_1[606] <= 0;lru_counter_2[606] <= 0;tag_1[606] <= 0;tag_2[606] <= 0;cache_mem_1[606] <= 0;cache_mem_2[606] <= 0;
    valid_1[607]  <=   0;valid_2[607]  <=   0;dirty_bit_1[607] <= 0;dirty_bit_2[607] <= 0;lru_counter_1[607] <= 0;lru_counter_2[607] <= 0;tag_1[607] <= 0;tag_2[607] <= 0;cache_mem_1[607] <= 0;cache_mem_2[607] <= 0;
    valid_1[608]  <=   0;valid_2[608]  <=   0;dirty_bit_1[608] <= 0;dirty_bit_2[608] <= 0;lru_counter_1[608] <= 0;lru_counter_2[608] <= 0;tag_1[608] <= 0;tag_2[608] <= 0;cache_mem_1[608] <= 0;cache_mem_2[608] <= 0;
    valid_1[609]  <=   0;valid_2[609]  <=   0;dirty_bit_1[609] <= 0;dirty_bit_2[609] <= 0;lru_counter_1[609] <= 0;lru_counter_2[609] <= 0;tag_1[609] <= 0;tag_2[609] <= 0;cache_mem_1[609] <= 0;cache_mem_2[609] <= 0;
    valid_1[610]  <=   0;valid_2[610]  <=   0;dirty_bit_1[610] <= 0;dirty_bit_2[610] <= 0;lru_counter_1[610] <= 0;lru_counter_2[610] <= 0;tag_1[610] <= 0;tag_2[610] <= 0;cache_mem_1[610] <= 0;cache_mem_2[610] <= 0;
    valid_1[611]  <=   0;valid_2[611]  <=   0;dirty_bit_1[611] <= 0;dirty_bit_2[611] <= 0;lru_counter_1[611] <= 0;lru_counter_2[611] <= 0;tag_1[611] <= 0;tag_2[611] <= 0;cache_mem_1[611] <= 0;cache_mem_2[611] <= 0;
    valid_1[612]  <=   0;valid_2[612]  <=   0;dirty_bit_1[612] <= 0;dirty_bit_2[612] <= 0;lru_counter_1[612] <= 0;lru_counter_2[612] <= 0;tag_1[612] <= 0;tag_2[612] <= 0;cache_mem_1[612] <= 0;cache_mem_2[612] <= 0;
    valid_1[613]  <=   0;valid_2[613]  <=   0;dirty_bit_1[613] <= 0;dirty_bit_2[613] <= 0;lru_counter_1[613] <= 0;lru_counter_2[613] <= 0;tag_1[613] <= 0;tag_2[613] <= 0;cache_mem_1[613] <= 0;cache_mem_2[613] <= 0;
    valid_1[614]  <=   0;valid_2[614]  <=   0;dirty_bit_1[614] <= 0;dirty_bit_2[614] <= 0;lru_counter_1[614] <= 0;lru_counter_2[614] <= 0;tag_1[614] <= 0;tag_2[614] <= 0;cache_mem_1[614] <= 0;cache_mem_2[614] <= 0;
    valid_1[615]  <=   0;valid_2[615]  <=   0;dirty_bit_1[615] <= 0;dirty_bit_2[615] <= 0;lru_counter_1[615] <= 0;lru_counter_2[615] <= 0;tag_1[615] <= 0;tag_2[615] <= 0;cache_mem_1[615] <= 0;cache_mem_2[615] <= 0;
    valid_1[616]  <=   0;valid_2[616]  <=   0;dirty_bit_1[616] <= 0;dirty_bit_2[616] <= 0;lru_counter_1[616] <= 0;lru_counter_2[616] <= 0;tag_1[616] <= 0;tag_2[616] <= 0;cache_mem_1[616] <= 0;cache_mem_2[616] <= 0;
    valid_1[617]  <=   0;valid_2[617]  <=   0;dirty_bit_1[617] <= 0;dirty_bit_2[617] <= 0;lru_counter_1[617] <= 0;lru_counter_2[617] <= 0;tag_1[617] <= 0;tag_2[617] <= 0;cache_mem_1[617] <= 0;cache_mem_2[617] <= 0;
    valid_1[618]  <=   0;valid_2[618]  <=   0;dirty_bit_1[618] <= 0;dirty_bit_2[618] <= 0;lru_counter_1[618] <= 0;lru_counter_2[618] <= 0;tag_1[618] <= 0;tag_2[618] <= 0;cache_mem_1[618] <= 0;cache_mem_2[618] <= 0;
    valid_1[619]  <=   0;valid_2[619]  <=   0;dirty_bit_1[619] <= 0;dirty_bit_2[619] <= 0;lru_counter_1[619] <= 0;lru_counter_2[619] <= 0;tag_1[619] <= 0;tag_2[619] <= 0;cache_mem_1[619] <= 0;cache_mem_2[619] <= 0;
    valid_1[620]  <=   0;valid_2[620]  <=   0;dirty_bit_1[620] <= 0;dirty_bit_2[620] <= 0;lru_counter_1[620] <= 0;lru_counter_2[620] <= 0;tag_1[620] <= 0;tag_2[620] <= 0;cache_mem_1[620] <= 0;cache_mem_2[620] <= 0;
    valid_1[621]  <=   0;valid_2[621]  <=   0;dirty_bit_1[621] <= 0;dirty_bit_2[621] <= 0;lru_counter_1[621] <= 0;lru_counter_2[621] <= 0;tag_1[621] <= 0;tag_2[621] <= 0;cache_mem_1[621] <= 0;cache_mem_2[621] <= 0;
    valid_1[622]  <=   0;valid_2[622]  <=   0;dirty_bit_1[622] <= 0;dirty_bit_2[622] <= 0;lru_counter_1[622] <= 0;lru_counter_2[622] <= 0;tag_1[622] <= 0;tag_2[622] <= 0;cache_mem_1[622] <= 0;cache_mem_2[622] <= 0;
    valid_1[623]  <=   0;valid_2[623]  <=   0;dirty_bit_1[623] <= 0;dirty_bit_2[623] <= 0;lru_counter_1[623] <= 0;lru_counter_2[623] <= 0;tag_1[623] <= 0;tag_2[623] <= 0;cache_mem_1[623] <= 0;cache_mem_2[623] <= 0;
    valid_1[624]  <=   0;valid_2[624]  <=   0;dirty_bit_1[624] <= 0;dirty_bit_2[624] <= 0;lru_counter_1[624] <= 0;lru_counter_2[624] <= 0;tag_1[624] <= 0;tag_2[624] <= 0;cache_mem_1[624] <= 0;cache_mem_2[624] <= 0;
    valid_1[625]  <=   0;valid_2[625]  <=   0;dirty_bit_1[625] <= 0;dirty_bit_2[625] <= 0;lru_counter_1[625] <= 0;lru_counter_2[625] <= 0;tag_1[625] <= 0;tag_2[625] <= 0;cache_mem_1[625] <= 0;cache_mem_2[625] <= 0;
    valid_1[626]  <=   0;valid_2[626]  <=   0;dirty_bit_1[626] <= 0;dirty_bit_2[626] <= 0;lru_counter_1[626] <= 0;lru_counter_2[626] <= 0;tag_1[626] <= 0;tag_2[626] <= 0;cache_mem_1[626] <= 0;cache_mem_2[626] <= 0;
    valid_1[627]  <=   0;valid_2[627]  <=   0;dirty_bit_1[627] <= 0;dirty_bit_2[627] <= 0;lru_counter_1[627] <= 0;lru_counter_2[627] <= 0;tag_1[627] <= 0;tag_2[627] <= 0;cache_mem_1[627] <= 0;cache_mem_2[627] <= 0;
    valid_1[628]  <=   0;valid_2[628]  <=   0;dirty_bit_1[628] <= 0;dirty_bit_2[628] <= 0;lru_counter_1[628] <= 0;lru_counter_2[628] <= 0;tag_1[628] <= 0;tag_2[628] <= 0;cache_mem_1[628] <= 0;cache_mem_2[628] <= 0;
    valid_1[629]  <=   0;valid_2[629]  <=   0;dirty_bit_1[629] <= 0;dirty_bit_2[629] <= 0;lru_counter_1[629] <= 0;lru_counter_2[629] <= 0;tag_1[629] <= 0;tag_2[629] <= 0;cache_mem_1[629] <= 0;cache_mem_2[629] <= 0;
    valid_1[630]  <=   0;valid_2[630]  <=   0;dirty_bit_1[630] <= 0;dirty_bit_2[630] <= 0;lru_counter_1[630] <= 0;lru_counter_2[630] <= 0;tag_1[630] <= 0;tag_2[630] <= 0;cache_mem_1[630] <= 0;cache_mem_2[630] <= 0;
    valid_1[631]  <=   0;valid_2[631]  <=   0;dirty_bit_1[631] <= 0;dirty_bit_2[631] <= 0;lru_counter_1[631] <= 0;lru_counter_2[631] <= 0;tag_1[631] <= 0;tag_2[631] <= 0;cache_mem_1[631] <= 0;cache_mem_2[631] <= 0;
    valid_1[632]  <=   0;valid_2[632]  <=   0;dirty_bit_1[632] <= 0;dirty_bit_2[632] <= 0;lru_counter_1[632] <= 0;lru_counter_2[632] <= 0;tag_1[632] <= 0;tag_2[632] <= 0;cache_mem_1[632] <= 0;cache_mem_2[632] <= 0;
    valid_1[633]  <=   0;valid_2[633]  <=   0;dirty_bit_1[633] <= 0;dirty_bit_2[633] <= 0;lru_counter_1[633] <= 0;lru_counter_2[633] <= 0;tag_1[633] <= 0;tag_2[633] <= 0;cache_mem_1[633] <= 0;cache_mem_2[633] <= 0;
    valid_1[634]  <=   0;valid_2[634]  <=   0;dirty_bit_1[634] <= 0;dirty_bit_2[634] <= 0;lru_counter_1[634] <= 0;lru_counter_2[634] <= 0;tag_1[634] <= 0;tag_2[634] <= 0;cache_mem_1[634] <= 0;cache_mem_2[634] <= 0;
    valid_1[635]  <=   0;valid_2[635]  <=   0;dirty_bit_1[635] <= 0;dirty_bit_2[635] <= 0;lru_counter_1[635] <= 0;lru_counter_2[635] <= 0;tag_1[635] <= 0;tag_2[635] <= 0;cache_mem_1[635] <= 0;cache_mem_2[635] <= 0;
    valid_1[636]  <=   0;valid_2[636]  <=   0;dirty_bit_1[636] <= 0;dirty_bit_2[636] <= 0;lru_counter_1[636] <= 0;lru_counter_2[636] <= 0;tag_1[636] <= 0;tag_2[636] <= 0;cache_mem_1[636] <= 0;cache_mem_2[636] <= 0;
    valid_1[637]  <=   0;valid_2[637]  <=   0;dirty_bit_1[637] <= 0;dirty_bit_2[637] <= 0;lru_counter_1[637] <= 0;lru_counter_2[637] <= 0;tag_1[637] <= 0;tag_2[637] <= 0;cache_mem_1[637] <= 0;cache_mem_2[637] <= 0;
    valid_1[638]  <=   0;valid_2[638]  <=   0;dirty_bit_1[638] <= 0;dirty_bit_2[638] <= 0;lru_counter_1[638] <= 0;lru_counter_2[638] <= 0;tag_1[638] <= 0;tag_2[638] <= 0;cache_mem_1[638] <= 0;cache_mem_2[638] <= 0;
    valid_1[639]  <=   0;valid_2[639]  <=   0;dirty_bit_1[639] <= 0;dirty_bit_2[639] <= 0;lru_counter_1[639] <= 0;lru_counter_2[639] <= 0;tag_1[639] <= 0;tag_2[639] <= 0;cache_mem_1[639] <= 0;cache_mem_2[639] <= 0;
    valid_1[640]  <=   0;valid_2[640]  <=   0;dirty_bit_1[640] <= 0;dirty_bit_2[640] <= 0;lru_counter_1[640] <= 0;lru_counter_2[640] <= 0;tag_1[640] <= 0;tag_2[640] <= 0;cache_mem_1[640] <= 0;cache_mem_2[640] <= 0;
    valid_1[641]  <=   0;valid_2[641]  <=   0;dirty_bit_1[641] <= 0;dirty_bit_2[641] <= 0;lru_counter_1[641] <= 0;lru_counter_2[641] <= 0;tag_1[641] <= 0;tag_2[641] <= 0;cache_mem_1[641] <= 0;cache_mem_2[641] <= 0;
    valid_1[642]  <=   0;valid_2[642]  <=   0;dirty_bit_1[642] <= 0;dirty_bit_2[642] <= 0;lru_counter_1[642] <= 0;lru_counter_2[642] <= 0;tag_1[642] <= 0;tag_2[642] <= 0;cache_mem_1[642] <= 0;cache_mem_2[642] <= 0;
    valid_1[643]  <=   0;valid_2[643]  <=   0;dirty_bit_1[643] <= 0;dirty_bit_2[643] <= 0;lru_counter_1[643] <= 0;lru_counter_2[643] <= 0;tag_1[643] <= 0;tag_2[643] <= 0;cache_mem_1[643] <= 0;cache_mem_2[643] <= 0;
    valid_1[644]  <=   0;valid_2[644]  <=   0;dirty_bit_1[644] <= 0;dirty_bit_2[644] <= 0;lru_counter_1[644] <= 0;lru_counter_2[644] <= 0;tag_1[644] <= 0;tag_2[644] <= 0;cache_mem_1[644] <= 0;cache_mem_2[644] <= 0;
    valid_1[645]  <=   0;valid_2[645]  <=   0;dirty_bit_1[645] <= 0;dirty_bit_2[645] <= 0;lru_counter_1[645] <= 0;lru_counter_2[645] <= 0;tag_1[645] <= 0;tag_2[645] <= 0;cache_mem_1[645] <= 0;cache_mem_2[645] <= 0;
    valid_1[646]  <=   0;valid_2[646]  <=   0;dirty_bit_1[646] <= 0;dirty_bit_2[646] <= 0;lru_counter_1[646] <= 0;lru_counter_2[646] <= 0;tag_1[646] <= 0;tag_2[646] <= 0;cache_mem_1[646] <= 0;cache_mem_2[646] <= 0;
    valid_1[647]  <=   0;valid_2[647]  <=   0;dirty_bit_1[647] <= 0;dirty_bit_2[647] <= 0;lru_counter_1[647] <= 0;lru_counter_2[647] <= 0;tag_1[647] <= 0;tag_2[647] <= 0;cache_mem_1[647] <= 0;cache_mem_2[647] <= 0;
    valid_1[648]  <=   0;valid_2[648]  <=   0;dirty_bit_1[648] <= 0;dirty_bit_2[648] <= 0;lru_counter_1[648] <= 0;lru_counter_2[648] <= 0;tag_1[648] <= 0;tag_2[648] <= 0;cache_mem_1[648] <= 0;cache_mem_2[648] <= 0;
    valid_1[649]  <=   0;valid_2[649]  <=   0;dirty_bit_1[649] <= 0;dirty_bit_2[649] <= 0;lru_counter_1[649] <= 0;lru_counter_2[649] <= 0;tag_1[649] <= 0;tag_2[649] <= 0;cache_mem_1[649] <= 0;cache_mem_2[649] <= 0;
    valid_1[650]  <=   0;valid_2[650]  <=   0;dirty_bit_1[650] <= 0;dirty_bit_2[650] <= 0;lru_counter_1[650] <= 0;lru_counter_2[650] <= 0;tag_1[650] <= 0;tag_2[650] <= 0;cache_mem_1[650] <= 0;cache_mem_2[650] <= 0;
    valid_1[651]  <=   0;valid_2[651]  <=   0;dirty_bit_1[651] <= 0;dirty_bit_2[651] <= 0;lru_counter_1[651] <= 0;lru_counter_2[651] <= 0;tag_1[651] <= 0;tag_2[651] <= 0;cache_mem_1[651] <= 0;cache_mem_2[651] <= 0;
    valid_1[652]  <=   0;valid_2[652]  <=   0;dirty_bit_1[652] <= 0;dirty_bit_2[652] <= 0;lru_counter_1[652] <= 0;lru_counter_2[652] <= 0;tag_1[652] <= 0;tag_2[652] <= 0;cache_mem_1[652] <= 0;cache_mem_2[652] <= 0;
    valid_1[653]  <=   0;valid_2[653]  <=   0;dirty_bit_1[653] <= 0;dirty_bit_2[653] <= 0;lru_counter_1[653] <= 0;lru_counter_2[653] <= 0;tag_1[653] <= 0;tag_2[653] <= 0;cache_mem_1[653] <= 0;cache_mem_2[653] <= 0;
    valid_1[654]  <=   0;valid_2[654]  <=   0;dirty_bit_1[654] <= 0;dirty_bit_2[654] <= 0;lru_counter_1[654] <= 0;lru_counter_2[654] <= 0;tag_1[654] <= 0;tag_2[654] <= 0;cache_mem_1[654] <= 0;cache_mem_2[654] <= 0;
    valid_1[655]  <=   0;valid_2[655]  <=   0;dirty_bit_1[655] <= 0;dirty_bit_2[655] <= 0;lru_counter_1[655] <= 0;lru_counter_2[655] <= 0;tag_1[655] <= 0;tag_2[655] <= 0;cache_mem_1[655] <= 0;cache_mem_2[655] <= 0;
    valid_1[656]  <=   0;valid_2[656]  <=   0;dirty_bit_1[656] <= 0;dirty_bit_2[656] <= 0;lru_counter_1[656] <= 0;lru_counter_2[656] <= 0;tag_1[656] <= 0;tag_2[656] <= 0;cache_mem_1[656] <= 0;cache_mem_2[656] <= 0;
    valid_1[657]  <=   0;valid_2[657]  <=   0;dirty_bit_1[657] <= 0;dirty_bit_2[657] <= 0;lru_counter_1[657] <= 0;lru_counter_2[657] <= 0;tag_1[657] <= 0;tag_2[657] <= 0;cache_mem_1[657] <= 0;cache_mem_2[657] <= 0;
    valid_1[658]  <=   0;valid_2[658]  <=   0;dirty_bit_1[658] <= 0;dirty_bit_2[658] <= 0;lru_counter_1[658] <= 0;lru_counter_2[658] <= 0;tag_1[658] <= 0;tag_2[658] <= 0;cache_mem_1[658] <= 0;cache_mem_2[658] <= 0;
    valid_1[659]  <=   0;valid_2[659]  <=   0;dirty_bit_1[659] <= 0;dirty_bit_2[659] <= 0;lru_counter_1[659] <= 0;lru_counter_2[659] <= 0;tag_1[659] <= 0;tag_2[659] <= 0;cache_mem_1[659] <= 0;cache_mem_2[659] <= 0;
    valid_1[660]  <=   0;valid_2[660]  <=   0;dirty_bit_1[660] <= 0;dirty_bit_2[660] <= 0;lru_counter_1[660] <= 0;lru_counter_2[660] <= 0;tag_1[660] <= 0;tag_2[660] <= 0;cache_mem_1[660] <= 0;cache_mem_2[660] <= 0;
    valid_1[661]  <=   0;valid_2[661]  <=   0;dirty_bit_1[661] <= 0;dirty_bit_2[661] <= 0;lru_counter_1[661] <= 0;lru_counter_2[661] <= 0;tag_1[661] <= 0;tag_2[661] <= 0;cache_mem_1[661] <= 0;cache_mem_2[661] <= 0;
    valid_1[662]  <=   0;valid_2[662]  <=   0;dirty_bit_1[662] <= 0;dirty_bit_2[662] <= 0;lru_counter_1[662] <= 0;lru_counter_2[662] <= 0;tag_1[662] <= 0;tag_2[662] <= 0;cache_mem_1[662] <= 0;cache_mem_2[662] <= 0;
    valid_1[663]  <=   0;valid_2[663]  <=   0;dirty_bit_1[663] <= 0;dirty_bit_2[663] <= 0;lru_counter_1[663] <= 0;lru_counter_2[663] <= 0;tag_1[663] <= 0;tag_2[663] <= 0;cache_mem_1[663] <= 0;cache_mem_2[663] <= 0;
    valid_1[664]  <=   0;valid_2[664]  <=   0;dirty_bit_1[664] <= 0;dirty_bit_2[664] <= 0;lru_counter_1[664] <= 0;lru_counter_2[664] <= 0;tag_1[664] <= 0;tag_2[664] <= 0;cache_mem_1[664] <= 0;cache_mem_2[664] <= 0;
    valid_1[665]  <=   0;valid_2[665]  <=   0;dirty_bit_1[665] <= 0;dirty_bit_2[665] <= 0;lru_counter_1[665] <= 0;lru_counter_2[665] <= 0;tag_1[665] <= 0;tag_2[665] <= 0;cache_mem_1[665] <= 0;cache_mem_2[665] <= 0;
    valid_1[666]  <=   0;valid_2[666]  <=   0;dirty_bit_1[666] <= 0;dirty_bit_2[666] <= 0;lru_counter_1[666] <= 0;lru_counter_2[666] <= 0;tag_1[666] <= 0;tag_2[666] <= 0;cache_mem_1[666] <= 0;cache_mem_2[666] <= 0;
    valid_1[667]  <=   0;valid_2[667]  <=   0;dirty_bit_1[667] <= 0;dirty_bit_2[667] <= 0;lru_counter_1[667] <= 0;lru_counter_2[667] <= 0;tag_1[667] <= 0;tag_2[667] <= 0;cache_mem_1[667] <= 0;cache_mem_2[667] <= 0;
    valid_1[668]  <=   0;valid_2[668]  <=   0;dirty_bit_1[668] <= 0;dirty_bit_2[668] <= 0;lru_counter_1[668] <= 0;lru_counter_2[668] <= 0;tag_1[668] <= 0;tag_2[668] <= 0;cache_mem_1[668] <= 0;cache_mem_2[668] <= 0;
    valid_1[669]  <=   0;valid_2[669]  <=   0;dirty_bit_1[669] <= 0;dirty_bit_2[669] <= 0;lru_counter_1[669] <= 0;lru_counter_2[669] <= 0;tag_1[669] <= 0;tag_2[669] <= 0;cache_mem_1[669] <= 0;cache_mem_2[669] <= 0;
    valid_1[670]  <=   0;valid_2[670]  <=   0;dirty_bit_1[670] <= 0;dirty_bit_2[670] <= 0;lru_counter_1[670] <= 0;lru_counter_2[670] <= 0;tag_1[670] <= 0;tag_2[670] <= 0;cache_mem_1[670] <= 0;cache_mem_2[670] <= 0;
    valid_1[671]  <=   0;valid_2[671]  <=   0;dirty_bit_1[671] <= 0;dirty_bit_2[671] <= 0;lru_counter_1[671] <= 0;lru_counter_2[671] <= 0;tag_1[671] <= 0;tag_2[671] <= 0;cache_mem_1[671] <= 0;cache_mem_2[671] <= 0;
    valid_1[672]  <=   0;valid_2[672]  <=   0;dirty_bit_1[672] <= 0;dirty_bit_2[672] <= 0;lru_counter_1[672] <= 0;lru_counter_2[672] <= 0;tag_1[672] <= 0;tag_2[672] <= 0;cache_mem_1[672] <= 0;cache_mem_2[672] <= 0;
    valid_1[673]  <=   0;valid_2[673]  <=   0;dirty_bit_1[673] <= 0;dirty_bit_2[673] <= 0;lru_counter_1[673] <= 0;lru_counter_2[673] <= 0;tag_1[673] <= 0;tag_2[673] <= 0;cache_mem_1[673] <= 0;cache_mem_2[673] <= 0;
    valid_1[674]  <=   0;valid_2[674]  <=   0;dirty_bit_1[674] <= 0;dirty_bit_2[674] <= 0;lru_counter_1[674] <= 0;lru_counter_2[674] <= 0;tag_1[674] <= 0;tag_2[674] <= 0;cache_mem_1[674] <= 0;cache_mem_2[674] <= 0;
    valid_1[675]  <=   0;valid_2[675]  <=   0;dirty_bit_1[675] <= 0;dirty_bit_2[675] <= 0;lru_counter_1[675] <= 0;lru_counter_2[675] <= 0;tag_1[675] <= 0;tag_2[675] <= 0;cache_mem_1[675] <= 0;cache_mem_2[675] <= 0;
    valid_1[676]  <=   0;valid_2[676]  <=   0;dirty_bit_1[676] <= 0;dirty_bit_2[676] <= 0;lru_counter_1[676] <= 0;lru_counter_2[676] <= 0;tag_1[676] <= 0;tag_2[676] <= 0;cache_mem_1[676] <= 0;cache_mem_2[676] <= 0;
    valid_1[677]  <=   0;valid_2[677]  <=   0;dirty_bit_1[677] <= 0;dirty_bit_2[677] <= 0;lru_counter_1[677] <= 0;lru_counter_2[677] <= 0;tag_1[677] <= 0;tag_2[677] <= 0;cache_mem_1[677] <= 0;cache_mem_2[677] <= 0;
    valid_1[678]  <=   0;valid_2[678]  <=   0;dirty_bit_1[678] <= 0;dirty_bit_2[678] <= 0;lru_counter_1[678] <= 0;lru_counter_2[678] <= 0;tag_1[678] <= 0;tag_2[678] <= 0;cache_mem_1[678] <= 0;cache_mem_2[678] <= 0;
    valid_1[679]  <=   0;valid_2[679]  <=   0;dirty_bit_1[679] <= 0;dirty_bit_2[679] <= 0;lru_counter_1[679] <= 0;lru_counter_2[679] <= 0;tag_1[679] <= 0;tag_2[679] <= 0;cache_mem_1[679] <= 0;cache_mem_2[679] <= 0;
    valid_1[680]  <=   0;valid_2[680]  <=   0;dirty_bit_1[680] <= 0;dirty_bit_2[680] <= 0;lru_counter_1[680] <= 0;lru_counter_2[680] <= 0;tag_1[680] <= 0;tag_2[680] <= 0;cache_mem_1[680] <= 0;cache_mem_2[680] <= 0;
    valid_1[681]  <=   0;valid_2[681]  <=   0;dirty_bit_1[681] <= 0;dirty_bit_2[681] <= 0;lru_counter_1[681] <= 0;lru_counter_2[681] <= 0;tag_1[681] <= 0;tag_2[681] <= 0;cache_mem_1[681] <= 0;cache_mem_2[681] <= 0;
    valid_1[682]  <=   0;valid_2[682]  <=   0;dirty_bit_1[682] <= 0;dirty_bit_2[682] <= 0;lru_counter_1[682] <= 0;lru_counter_2[682] <= 0;tag_1[682] <= 0;tag_2[682] <= 0;cache_mem_1[682] <= 0;cache_mem_2[682] <= 0;
    valid_1[683]  <=   0;valid_2[683]  <=   0;dirty_bit_1[683] <= 0;dirty_bit_2[683] <= 0;lru_counter_1[683] <= 0;lru_counter_2[683] <= 0;tag_1[683] <= 0;tag_2[683] <= 0;cache_mem_1[683] <= 0;cache_mem_2[683] <= 0;
    valid_1[684]  <=   0;valid_2[684]  <=   0;dirty_bit_1[684] <= 0;dirty_bit_2[684] <= 0;lru_counter_1[684] <= 0;lru_counter_2[684] <= 0;tag_1[684] <= 0;tag_2[684] <= 0;cache_mem_1[684] <= 0;cache_mem_2[684] <= 0;
    valid_1[685]  <=   0;valid_2[685]  <=   0;dirty_bit_1[685] <= 0;dirty_bit_2[685] <= 0;lru_counter_1[685] <= 0;lru_counter_2[685] <= 0;tag_1[685] <= 0;tag_2[685] <= 0;cache_mem_1[685] <= 0;cache_mem_2[685] <= 0;
    valid_1[686]  <=   0;valid_2[686]  <=   0;dirty_bit_1[686] <= 0;dirty_bit_2[686] <= 0;lru_counter_1[686] <= 0;lru_counter_2[686] <= 0;tag_1[686] <= 0;tag_2[686] <= 0;cache_mem_1[686] <= 0;cache_mem_2[686] <= 0;
    valid_1[687]  <=   0;valid_2[687]  <=   0;dirty_bit_1[687] <= 0;dirty_bit_2[687] <= 0;lru_counter_1[687] <= 0;lru_counter_2[687] <= 0;tag_1[687] <= 0;tag_2[687] <= 0;cache_mem_1[687] <= 0;cache_mem_2[687] <= 0;
    valid_1[688]  <=   0;valid_2[688]  <=   0;dirty_bit_1[688] <= 0;dirty_bit_2[688] <= 0;lru_counter_1[688] <= 0;lru_counter_2[688] <= 0;tag_1[688] <= 0;tag_2[688] <= 0;cache_mem_1[688] <= 0;cache_mem_2[688] <= 0;
    valid_1[689]  <=   0;valid_2[689]  <=   0;dirty_bit_1[689] <= 0;dirty_bit_2[689] <= 0;lru_counter_1[689] <= 0;lru_counter_2[689] <= 0;tag_1[689] <= 0;tag_2[689] <= 0;cache_mem_1[689] <= 0;cache_mem_2[689] <= 0;
    valid_1[690]  <=   0;valid_2[690]  <=   0;dirty_bit_1[690] <= 0;dirty_bit_2[690] <= 0;lru_counter_1[690] <= 0;lru_counter_2[690] <= 0;tag_1[690] <= 0;tag_2[690] <= 0;cache_mem_1[690] <= 0;cache_mem_2[690] <= 0;
    valid_1[691]  <=   0;valid_2[691]  <=   0;dirty_bit_1[691] <= 0;dirty_bit_2[691] <= 0;lru_counter_1[691] <= 0;lru_counter_2[691] <= 0;tag_1[691] <= 0;tag_2[691] <= 0;cache_mem_1[691] <= 0;cache_mem_2[691] <= 0;
    valid_1[692]  <=   0;valid_2[692]  <=   0;dirty_bit_1[692] <= 0;dirty_bit_2[692] <= 0;lru_counter_1[692] <= 0;lru_counter_2[692] <= 0;tag_1[692] <= 0;tag_2[692] <= 0;cache_mem_1[692] <= 0;cache_mem_2[692] <= 0;
    valid_1[693]  <=   0;valid_2[693]  <=   0;dirty_bit_1[693] <= 0;dirty_bit_2[693] <= 0;lru_counter_1[693] <= 0;lru_counter_2[693] <= 0;tag_1[693] <= 0;tag_2[693] <= 0;cache_mem_1[693] <= 0;cache_mem_2[693] <= 0;
    valid_1[694]  <=   0;valid_2[694]  <=   0;dirty_bit_1[694] <= 0;dirty_bit_2[694] <= 0;lru_counter_1[694] <= 0;lru_counter_2[694] <= 0;tag_1[694] <= 0;tag_2[694] <= 0;cache_mem_1[694] <= 0;cache_mem_2[694] <= 0;
    valid_1[695]  <=   0;valid_2[695]  <=   0;dirty_bit_1[695] <= 0;dirty_bit_2[695] <= 0;lru_counter_1[695] <= 0;lru_counter_2[695] <= 0;tag_1[695] <= 0;tag_2[695] <= 0;cache_mem_1[695] <= 0;cache_mem_2[695] <= 0;
    valid_1[696]  <=   0;valid_2[696]  <=   0;dirty_bit_1[696] <= 0;dirty_bit_2[696] <= 0;lru_counter_1[696] <= 0;lru_counter_2[696] <= 0;tag_1[696] <= 0;tag_2[696] <= 0;cache_mem_1[696] <= 0;cache_mem_2[696] <= 0;
    valid_1[697]  <=   0;valid_2[697]  <=   0;dirty_bit_1[697] <= 0;dirty_bit_2[697] <= 0;lru_counter_1[697] <= 0;lru_counter_2[697] <= 0;tag_1[697] <= 0;tag_2[697] <= 0;cache_mem_1[697] <= 0;cache_mem_2[697] <= 0;
    valid_1[698]  <=   0;valid_2[698]  <=   0;dirty_bit_1[698] <= 0;dirty_bit_2[698] <= 0;lru_counter_1[698] <= 0;lru_counter_2[698] <= 0;tag_1[698] <= 0;tag_2[698] <= 0;cache_mem_1[698] <= 0;cache_mem_2[698] <= 0;
    valid_1[699]  <=   0;valid_2[699]  <=   0;dirty_bit_1[699] <= 0;dirty_bit_2[699] <= 0;lru_counter_1[699] <= 0;lru_counter_2[699] <= 0;tag_1[699] <= 0;tag_2[699] <= 0;cache_mem_1[699] <= 0;cache_mem_2[699] <= 0;
    valid_1[700]  <=   0;valid_2[700]  <=   0;dirty_bit_1[700] <= 0;dirty_bit_2[700] <= 0;lru_counter_1[700] <= 0;lru_counter_2[700] <= 0;tag_1[700] <= 0;tag_2[700] <= 0;cache_mem_1[700] <= 0;cache_mem_2[700] <= 0;
    valid_1[701]  <=   0;valid_2[701]  <=   0;dirty_bit_1[701] <= 0;dirty_bit_2[701] <= 0;lru_counter_1[701] <= 0;lru_counter_2[701] <= 0;tag_1[701] <= 0;tag_2[701] <= 0;cache_mem_1[701] <= 0;cache_mem_2[701] <= 0;
    valid_1[702]  <=   0;valid_2[702]  <=   0;dirty_bit_1[702] <= 0;dirty_bit_2[702] <= 0;lru_counter_1[702] <= 0;lru_counter_2[702] <= 0;tag_1[702] <= 0;tag_2[702] <= 0;cache_mem_1[702] <= 0;cache_mem_2[702] <= 0;
    valid_1[703]  <=   0;valid_2[703]  <=   0;dirty_bit_1[703] <= 0;dirty_bit_2[703] <= 0;lru_counter_1[703] <= 0;lru_counter_2[703] <= 0;tag_1[703] <= 0;tag_2[703] <= 0;cache_mem_1[703] <= 0;cache_mem_2[703] <= 0;
    valid_1[704]  <=   0;valid_2[704]  <=   0;dirty_bit_1[704] <= 0;dirty_bit_2[704] <= 0;lru_counter_1[704] <= 0;lru_counter_2[704] <= 0;tag_1[704] <= 0;tag_2[704] <= 0;cache_mem_1[704] <= 0;cache_mem_2[704] <= 0;
    valid_1[705]  <=   0;valid_2[705]  <=   0;dirty_bit_1[705] <= 0;dirty_bit_2[705] <= 0;lru_counter_1[705] <= 0;lru_counter_2[705] <= 0;tag_1[705] <= 0;tag_2[705] <= 0;cache_mem_1[705] <= 0;cache_mem_2[705] <= 0;
    valid_1[706]  <=   0;valid_2[706]  <=   0;dirty_bit_1[706] <= 0;dirty_bit_2[706] <= 0;lru_counter_1[706] <= 0;lru_counter_2[706] <= 0;tag_1[706] <= 0;tag_2[706] <= 0;cache_mem_1[706] <= 0;cache_mem_2[706] <= 0;
    valid_1[707]  <=   0;valid_2[707]  <=   0;dirty_bit_1[707] <= 0;dirty_bit_2[707] <= 0;lru_counter_1[707] <= 0;lru_counter_2[707] <= 0;tag_1[707] <= 0;tag_2[707] <= 0;cache_mem_1[707] <= 0;cache_mem_2[707] <= 0;
    valid_1[708]  <=   0;valid_2[708]  <=   0;dirty_bit_1[708] <= 0;dirty_bit_2[708] <= 0;lru_counter_1[708] <= 0;lru_counter_2[708] <= 0;tag_1[708] <= 0;tag_2[708] <= 0;cache_mem_1[708] <= 0;cache_mem_2[708] <= 0;
    valid_1[709]  <=   0;valid_2[709]  <=   0;dirty_bit_1[709] <= 0;dirty_bit_2[709] <= 0;lru_counter_1[709] <= 0;lru_counter_2[709] <= 0;tag_1[709] <= 0;tag_2[709] <= 0;cache_mem_1[709] <= 0;cache_mem_2[709] <= 0;
    valid_1[710]  <=   0;valid_2[710]  <=   0;dirty_bit_1[710] <= 0;dirty_bit_2[710] <= 0;lru_counter_1[710] <= 0;lru_counter_2[710] <= 0;tag_1[710] <= 0;tag_2[710] <= 0;cache_mem_1[710] <= 0;cache_mem_2[710] <= 0;
    valid_1[711]  <=   0;valid_2[711]  <=   0;dirty_bit_1[711] <= 0;dirty_bit_2[711] <= 0;lru_counter_1[711] <= 0;lru_counter_2[711] <= 0;tag_1[711] <= 0;tag_2[711] <= 0;cache_mem_1[711] <= 0;cache_mem_2[711] <= 0;
    valid_1[712]  <=   0;valid_2[712]  <=   0;dirty_bit_1[712] <= 0;dirty_bit_2[712] <= 0;lru_counter_1[712] <= 0;lru_counter_2[712] <= 0;tag_1[712] <= 0;tag_2[712] <= 0;cache_mem_1[712] <= 0;cache_mem_2[712] <= 0;
    valid_1[713]  <=   0;valid_2[713]  <=   0;dirty_bit_1[713] <= 0;dirty_bit_2[713] <= 0;lru_counter_1[713] <= 0;lru_counter_2[713] <= 0;tag_1[713] <= 0;tag_2[713] <= 0;cache_mem_1[713] <= 0;cache_mem_2[713] <= 0;
    valid_1[714]  <=   0;valid_2[714]  <=   0;dirty_bit_1[714] <= 0;dirty_bit_2[714] <= 0;lru_counter_1[714] <= 0;lru_counter_2[714] <= 0;tag_1[714] <= 0;tag_2[714] <= 0;cache_mem_1[714] <= 0;cache_mem_2[714] <= 0;
    valid_1[715]  <=   0;valid_2[715]  <=   0;dirty_bit_1[715] <= 0;dirty_bit_2[715] <= 0;lru_counter_1[715] <= 0;lru_counter_2[715] <= 0;tag_1[715] <= 0;tag_2[715] <= 0;cache_mem_1[715] <= 0;cache_mem_2[715] <= 0;
    valid_1[716]  <=   0;valid_2[716]  <=   0;dirty_bit_1[716] <= 0;dirty_bit_2[716] <= 0;lru_counter_1[716] <= 0;lru_counter_2[716] <= 0;tag_1[716] <= 0;tag_2[716] <= 0;cache_mem_1[716] <= 0;cache_mem_2[716] <= 0;
    valid_1[717]  <=   0;valid_2[717]  <=   0;dirty_bit_1[717] <= 0;dirty_bit_2[717] <= 0;lru_counter_1[717] <= 0;lru_counter_2[717] <= 0;tag_1[717] <= 0;tag_2[717] <= 0;cache_mem_1[717] <= 0;cache_mem_2[717] <= 0;
    valid_1[718]  <=   0;valid_2[718]  <=   0;dirty_bit_1[718] <= 0;dirty_bit_2[718] <= 0;lru_counter_1[718] <= 0;lru_counter_2[718] <= 0;tag_1[718] <= 0;tag_2[718] <= 0;cache_mem_1[718] <= 0;cache_mem_2[718] <= 0;
    valid_1[719]  <=   0;valid_2[719]  <=   0;dirty_bit_1[719] <= 0;dirty_bit_2[719] <= 0;lru_counter_1[719] <= 0;lru_counter_2[719] <= 0;tag_1[719] <= 0;tag_2[719] <= 0;cache_mem_1[719] <= 0;cache_mem_2[719] <= 0;
    valid_1[720]  <=   0;valid_2[720]  <=   0;dirty_bit_1[720] <= 0;dirty_bit_2[720] <= 0;lru_counter_1[720] <= 0;lru_counter_2[720] <= 0;tag_1[720] <= 0;tag_2[720] <= 0;cache_mem_1[720] <= 0;cache_mem_2[720] <= 0;
    valid_1[721]  <=   0;valid_2[721]  <=   0;dirty_bit_1[721] <= 0;dirty_bit_2[721] <= 0;lru_counter_1[721] <= 0;lru_counter_2[721] <= 0;tag_1[721] <= 0;tag_2[721] <= 0;cache_mem_1[721] <= 0;cache_mem_2[721] <= 0;
    valid_1[722]  <=   0;valid_2[722]  <=   0;dirty_bit_1[722] <= 0;dirty_bit_2[722] <= 0;lru_counter_1[722] <= 0;lru_counter_2[722] <= 0;tag_1[722] <= 0;tag_2[722] <= 0;cache_mem_1[722] <= 0;cache_mem_2[722] <= 0;
    valid_1[723]  <=   0;valid_2[723]  <=   0;dirty_bit_1[723] <= 0;dirty_bit_2[723] <= 0;lru_counter_1[723] <= 0;lru_counter_2[723] <= 0;tag_1[723] <= 0;tag_2[723] <= 0;cache_mem_1[723] <= 0;cache_mem_2[723] <= 0;
    valid_1[724]  <=   0;valid_2[724]  <=   0;dirty_bit_1[724] <= 0;dirty_bit_2[724] <= 0;lru_counter_1[724] <= 0;lru_counter_2[724] <= 0;tag_1[724] <= 0;tag_2[724] <= 0;cache_mem_1[724] <= 0;cache_mem_2[724] <= 0;
    valid_1[725]  <=   0;valid_2[725]  <=   0;dirty_bit_1[725] <= 0;dirty_bit_2[725] <= 0;lru_counter_1[725] <= 0;lru_counter_2[725] <= 0;tag_1[725] <= 0;tag_2[725] <= 0;cache_mem_1[725] <= 0;cache_mem_2[725] <= 0;
    valid_1[726]  <=   0;valid_2[726]  <=   0;dirty_bit_1[726] <= 0;dirty_bit_2[726] <= 0;lru_counter_1[726] <= 0;lru_counter_2[726] <= 0;tag_1[726] <= 0;tag_2[726] <= 0;cache_mem_1[726] <= 0;cache_mem_2[726] <= 0;
    valid_1[727]  <=   0;valid_2[727]  <=   0;dirty_bit_1[727] <= 0;dirty_bit_2[727] <= 0;lru_counter_1[727] <= 0;lru_counter_2[727] <= 0;tag_1[727] <= 0;tag_2[727] <= 0;cache_mem_1[727] <= 0;cache_mem_2[727] <= 0;
    valid_1[728]  <=   0;valid_2[728]  <=   0;dirty_bit_1[728] <= 0;dirty_bit_2[728] <= 0;lru_counter_1[728] <= 0;lru_counter_2[728] <= 0;tag_1[728] <= 0;tag_2[728] <= 0;cache_mem_1[728] <= 0;cache_mem_2[728] <= 0;
    valid_1[729]  <=   0;valid_2[729]  <=   0;dirty_bit_1[729] <= 0;dirty_bit_2[729] <= 0;lru_counter_1[729] <= 0;lru_counter_2[729] <= 0;tag_1[729] <= 0;tag_2[729] <= 0;cache_mem_1[729] <= 0;cache_mem_2[729] <= 0;
    valid_1[730]  <=   0;valid_2[730]  <=   0;dirty_bit_1[730] <= 0;dirty_bit_2[730] <= 0;lru_counter_1[730] <= 0;lru_counter_2[730] <= 0;tag_1[730] <= 0;tag_2[730] <= 0;cache_mem_1[730] <= 0;cache_mem_2[730] <= 0;
    valid_1[731]  <=   0;valid_2[731]  <=   0;dirty_bit_1[731] <= 0;dirty_bit_2[731] <= 0;lru_counter_1[731] <= 0;lru_counter_2[731] <= 0;tag_1[731] <= 0;tag_2[731] <= 0;cache_mem_1[731] <= 0;cache_mem_2[731] <= 0;
    valid_1[732]  <=   0;valid_2[732]  <=   0;dirty_bit_1[732] <= 0;dirty_bit_2[732] <= 0;lru_counter_1[732] <= 0;lru_counter_2[732] <= 0;tag_1[732] <= 0;tag_2[732] <= 0;cache_mem_1[732] <= 0;cache_mem_2[732] <= 0;
    valid_1[733]  <=   0;valid_2[733]  <=   0;dirty_bit_1[733] <= 0;dirty_bit_2[733] <= 0;lru_counter_1[733] <= 0;lru_counter_2[733] <= 0;tag_1[733] <= 0;tag_2[733] <= 0;cache_mem_1[733] <= 0;cache_mem_2[733] <= 0;
    valid_1[734]  <=   0;valid_2[734]  <=   0;dirty_bit_1[734] <= 0;dirty_bit_2[734] <= 0;lru_counter_1[734] <= 0;lru_counter_2[734] <= 0;tag_1[734] <= 0;tag_2[734] <= 0;cache_mem_1[734] <= 0;cache_mem_2[734] <= 0;
    valid_1[735]  <=   0;valid_2[735]  <=   0;dirty_bit_1[735] <= 0;dirty_bit_2[735] <= 0;lru_counter_1[735] <= 0;lru_counter_2[735] <= 0;tag_1[735] <= 0;tag_2[735] <= 0;cache_mem_1[735] <= 0;cache_mem_2[735] <= 0;
    valid_1[736]  <=   0;valid_2[736]  <=   0;dirty_bit_1[736] <= 0;dirty_bit_2[736] <= 0;lru_counter_1[736] <= 0;lru_counter_2[736] <= 0;tag_1[736] <= 0;tag_2[736] <= 0;cache_mem_1[736] <= 0;cache_mem_2[736] <= 0;
    valid_1[737]  <=   0;valid_2[737]  <=   0;dirty_bit_1[737] <= 0;dirty_bit_2[737] <= 0;lru_counter_1[737] <= 0;lru_counter_2[737] <= 0;tag_1[737] <= 0;tag_2[737] <= 0;cache_mem_1[737] <= 0;cache_mem_2[737] <= 0;
    valid_1[738]  <=   0;valid_2[738]  <=   0;dirty_bit_1[738] <= 0;dirty_bit_2[738] <= 0;lru_counter_1[738] <= 0;lru_counter_2[738] <= 0;tag_1[738] <= 0;tag_2[738] <= 0;cache_mem_1[738] <= 0;cache_mem_2[738] <= 0;
    valid_1[739]  <=   0;valid_2[739]  <=   0;dirty_bit_1[739] <= 0;dirty_bit_2[739] <= 0;lru_counter_1[739] <= 0;lru_counter_2[739] <= 0;tag_1[739] <= 0;tag_2[739] <= 0;cache_mem_1[739] <= 0;cache_mem_2[739] <= 0;
    valid_1[740]  <=   0;valid_2[740]  <=   0;dirty_bit_1[740] <= 0;dirty_bit_2[740] <= 0;lru_counter_1[740] <= 0;lru_counter_2[740] <= 0;tag_1[740] <= 0;tag_2[740] <= 0;cache_mem_1[740] <= 0;cache_mem_2[740] <= 0;
    valid_1[741]  <=   0;valid_2[741]  <=   0;dirty_bit_1[741] <= 0;dirty_bit_2[741] <= 0;lru_counter_1[741] <= 0;lru_counter_2[741] <= 0;tag_1[741] <= 0;tag_2[741] <= 0;cache_mem_1[741] <= 0;cache_mem_2[741] <= 0;
    valid_1[742]  <=   0;valid_2[742]  <=   0;dirty_bit_1[742] <= 0;dirty_bit_2[742] <= 0;lru_counter_1[742] <= 0;lru_counter_2[742] <= 0;tag_1[742] <= 0;tag_2[742] <= 0;cache_mem_1[742] <= 0;cache_mem_2[742] <= 0;
    valid_1[743]  <=   0;valid_2[743]  <=   0;dirty_bit_1[743] <= 0;dirty_bit_2[743] <= 0;lru_counter_1[743] <= 0;lru_counter_2[743] <= 0;tag_1[743] <= 0;tag_2[743] <= 0;cache_mem_1[743] <= 0;cache_mem_2[743] <= 0;
    valid_1[744]  <=   0;valid_2[744]  <=   0;dirty_bit_1[744] <= 0;dirty_bit_2[744] <= 0;lru_counter_1[744] <= 0;lru_counter_2[744] <= 0;tag_1[744] <= 0;tag_2[744] <= 0;cache_mem_1[744] <= 0;cache_mem_2[744] <= 0;
    valid_1[745]  <=   0;valid_2[745]  <=   0;dirty_bit_1[745] <= 0;dirty_bit_2[745] <= 0;lru_counter_1[745] <= 0;lru_counter_2[745] <= 0;tag_1[745] <= 0;tag_2[745] <= 0;cache_mem_1[745] <= 0;cache_mem_2[745] <= 0;
    valid_1[746]  <=   0;valid_2[746]  <=   0;dirty_bit_1[746] <= 0;dirty_bit_2[746] <= 0;lru_counter_1[746] <= 0;lru_counter_2[746] <= 0;tag_1[746] <= 0;tag_2[746] <= 0;cache_mem_1[746] <= 0;cache_mem_2[746] <= 0;
    valid_1[747]  <=   0;valid_2[747]  <=   0;dirty_bit_1[747] <= 0;dirty_bit_2[747] <= 0;lru_counter_1[747] <= 0;lru_counter_2[747] <= 0;tag_1[747] <= 0;tag_2[747] <= 0;cache_mem_1[747] <= 0;cache_mem_2[747] <= 0;
    valid_1[748]  <=   0;valid_2[748]  <=   0;dirty_bit_1[748] <= 0;dirty_bit_2[748] <= 0;lru_counter_1[748] <= 0;lru_counter_2[748] <= 0;tag_1[748] <= 0;tag_2[748] <= 0;cache_mem_1[748] <= 0;cache_mem_2[748] <= 0;
    valid_1[749]  <=   0;valid_2[749]  <=   0;dirty_bit_1[749] <= 0;dirty_bit_2[749] <= 0;lru_counter_1[749] <= 0;lru_counter_2[749] <= 0;tag_1[749] <= 0;tag_2[749] <= 0;cache_mem_1[749] <= 0;cache_mem_2[749] <= 0;
    valid_1[750]  <=   0;valid_2[750]  <=   0;dirty_bit_1[750] <= 0;dirty_bit_2[750] <= 0;lru_counter_1[750] <= 0;lru_counter_2[750] <= 0;tag_1[750] <= 0;tag_2[750] <= 0;cache_mem_1[750] <= 0;cache_mem_2[750] <= 0;
    valid_1[751]  <=   0;valid_2[751]  <=   0;dirty_bit_1[751] <= 0;dirty_bit_2[751] <= 0;lru_counter_1[751] <= 0;lru_counter_2[751] <= 0;tag_1[751] <= 0;tag_2[751] <= 0;cache_mem_1[751] <= 0;cache_mem_2[751] <= 0;
    valid_1[752]  <=   0;valid_2[752]  <=   0;dirty_bit_1[752] <= 0;dirty_bit_2[752] <= 0;lru_counter_1[752] <= 0;lru_counter_2[752] <= 0;tag_1[752] <= 0;tag_2[752] <= 0;cache_mem_1[752] <= 0;cache_mem_2[752] <= 0;
    valid_1[753]  <=   0;valid_2[753]  <=   0;dirty_bit_1[753] <= 0;dirty_bit_2[753] <= 0;lru_counter_1[753] <= 0;lru_counter_2[753] <= 0;tag_1[753] <= 0;tag_2[753] <= 0;cache_mem_1[753] <= 0;cache_mem_2[753] <= 0;
    valid_1[754]  <=   0;valid_2[754]  <=   0;dirty_bit_1[754] <= 0;dirty_bit_2[754] <= 0;lru_counter_1[754] <= 0;lru_counter_2[754] <= 0;tag_1[754] <= 0;tag_2[754] <= 0;cache_mem_1[754] <= 0;cache_mem_2[754] <= 0;
    valid_1[755]  <=   0;valid_2[755]  <=   0;dirty_bit_1[755] <= 0;dirty_bit_2[755] <= 0;lru_counter_1[755] <= 0;lru_counter_2[755] <= 0;tag_1[755] <= 0;tag_2[755] <= 0;cache_mem_1[755] <= 0;cache_mem_2[755] <= 0;
    valid_1[756]  <=   0;valid_2[756]  <=   0;dirty_bit_1[756] <= 0;dirty_bit_2[756] <= 0;lru_counter_1[756] <= 0;lru_counter_2[756] <= 0;tag_1[756] <= 0;tag_2[756] <= 0;cache_mem_1[756] <= 0;cache_mem_2[756] <= 0;
    valid_1[757]  <=   0;valid_2[757]  <=   0;dirty_bit_1[757] <= 0;dirty_bit_2[757] <= 0;lru_counter_1[757] <= 0;lru_counter_2[757] <= 0;tag_1[757] <= 0;tag_2[757] <= 0;cache_mem_1[757] <= 0;cache_mem_2[757] <= 0;
    valid_1[758]  <=   0;valid_2[758]  <=   0;dirty_bit_1[758] <= 0;dirty_bit_2[758] <= 0;lru_counter_1[758] <= 0;lru_counter_2[758] <= 0;tag_1[758] <= 0;tag_2[758] <= 0;cache_mem_1[758] <= 0;cache_mem_2[758] <= 0;
    valid_1[759]  <=   0;valid_2[759]  <=   0;dirty_bit_1[759] <= 0;dirty_bit_2[759] <= 0;lru_counter_1[759] <= 0;lru_counter_2[759] <= 0;tag_1[759] <= 0;tag_2[759] <= 0;cache_mem_1[759] <= 0;cache_mem_2[759] <= 0;
    valid_1[760]  <=   0;valid_2[760]  <=   0;dirty_bit_1[760] <= 0;dirty_bit_2[760] <= 0;lru_counter_1[760] <= 0;lru_counter_2[760] <= 0;tag_1[760] <= 0;tag_2[760] <= 0;cache_mem_1[760] <= 0;cache_mem_2[760] <= 0;
    valid_1[761]  <=   0;valid_2[761]  <=   0;dirty_bit_1[761] <= 0;dirty_bit_2[761] <= 0;lru_counter_1[761] <= 0;lru_counter_2[761] <= 0;tag_1[761] <= 0;tag_2[761] <= 0;cache_mem_1[761] <= 0;cache_mem_2[761] <= 0;
    valid_1[762]  <=   0;valid_2[762]  <=   0;dirty_bit_1[762] <= 0;dirty_bit_2[762] <= 0;lru_counter_1[762] <= 0;lru_counter_2[762] <= 0;tag_1[762] <= 0;tag_2[762] <= 0;cache_mem_1[762] <= 0;cache_mem_2[762] <= 0;
    valid_1[763]  <=   0;valid_2[763]  <=   0;dirty_bit_1[763] <= 0;dirty_bit_2[763] <= 0;lru_counter_1[763] <= 0;lru_counter_2[763] <= 0;tag_1[763] <= 0;tag_2[763] <= 0;cache_mem_1[763] <= 0;cache_mem_2[763] <= 0;
    valid_1[764]  <=   0;valid_2[764]  <=   0;dirty_bit_1[764] <= 0;dirty_bit_2[764] <= 0;lru_counter_1[764] <= 0;lru_counter_2[764] <= 0;tag_1[764] <= 0;tag_2[764] <= 0;cache_mem_1[764] <= 0;cache_mem_2[764] <= 0;
    valid_1[765]  <=   0;valid_2[765]  <=   0;dirty_bit_1[765] <= 0;dirty_bit_2[765] <= 0;lru_counter_1[765] <= 0;lru_counter_2[765] <= 0;tag_1[765] <= 0;tag_2[765] <= 0;cache_mem_1[765] <= 0;cache_mem_2[765] <= 0;
    valid_1[766]  <=   0;valid_2[766]  <=   0;dirty_bit_1[766] <= 0;dirty_bit_2[766] <= 0;lru_counter_1[766] <= 0;lru_counter_2[766] <= 0;tag_1[766] <= 0;tag_2[766] <= 0;cache_mem_1[766] <= 0;cache_mem_2[766] <= 0;
    valid_1[767]  <=   0;valid_2[767]  <=   0;dirty_bit_1[767] <= 0;dirty_bit_2[767] <= 0;lru_counter_1[767] <= 0;lru_counter_2[767] <= 0;tag_1[767] <= 0;tag_2[767] <= 0;cache_mem_1[767] <= 0;cache_mem_2[767] <= 0;
    valid_1[768]  <=   0;valid_2[768]  <=   0;dirty_bit_1[768] <= 0;dirty_bit_2[768] <= 0;lru_counter_1[768] <= 0;lru_counter_2[768] <= 0;tag_1[768] <= 0;tag_2[768] <= 0;cache_mem_1[768] <= 0;cache_mem_2[768] <= 0;
    valid_1[769]  <=   0;valid_2[769]  <=   0;dirty_bit_1[769] <= 0;dirty_bit_2[769] <= 0;lru_counter_1[769] <= 0;lru_counter_2[769] <= 0;tag_1[769] <= 0;tag_2[769] <= 0;cache_mem_1[769] <= 0;cache_mem_2[769] <= 0;
    valid_1[770]  <=   0;valid_2[770]  <=   0;dirty_bit_1[770] <= 0;dirty_bit_2[770] <= 0;lru_counter_1[770] <= 0;lru_counter_2[770] <= 0;tag_1[770] <= 0;tag_2[770] <= 0;cache_mem_1[770] <= 0;cache_mem_2[770] <= 0;
    valid_1[771]  <=   0;valid_2[771]  <=   0;dirty_bit_1[771] <= 0;dirty_bit_2[771] <= 0;lru_counter_1[771] <= 0;lru_counter_2[771] <= 0;tag_1[771] <= 0;tag_2[771] <= 0;cache_mem_1[771] <= 0;cache_mem_2[771] <= 0;
    valid_1[772]  <=   0;valid_2[772]  <=   0;dirty_bit_1[772] <= 0;dirty_bit_2[772] <= 0;lru_counter_1[772] <= 0;lru_counter_2[772] <= 0;tag_1[772] <= 0;tag_2[772] <= 0;cache_mem_1[772] <= 0;cache_mem_2[772] <= 0;
    valid_1[773]  <=   0;valid_2[773]  <=   0;dirty_bit_1[773] <= 0;dirty_bit_2[773] <= 0;lru_counter_1[773] <= 0;lru_counter_2[773] <= 0;tag_1[773] <= 0;tag_2[773] <= 0;cache_mem_1[773] <= 0;cache_mem_2[773] <= 0;
    valid_1[774]  <=   0;valid_2[774]  <=   0;dirty_bit_1[774] <= 0;dirty_bit_2[774] <= 0;lru_counter_1[774] <= 0;lru_counter_2[774] <= 0;tag_1[774] <= 0;tag_2[774] <= 0;cache_mem_1[774] <= 0;cache_mem_2[774] <= 0;
    valid_1[775]  <=   0;valid_2[775]  <=   0;dirty_bit_1[775] <= 0;dirty_bit_2[775] <= 0;lru_counter_1[775] <= 0;lru_counter_2[775] <= 0;tag_1[775] <= 0;tag_2[775] <= 0;cache_mem_1[775] <= 0;cache_mem_2[775] <= 0;
    valid_1[776]  <=   0;valid_2[776]  <=   0;dirty_bit_1[776] <= 0;dirty_bit_2[776] <= 0;lru_counter_1[776] <= 0;lru_counter_2[776] <= 0;tag_1[776] <= 0;tag_2[776] <= 0;cache_mem_1[776] <= 0;cache_mem_2[776] <= 0;
    valid_1[777]  <=   0;valid_2[777]  <=   0;dirty_bit_1[777] <= 0;dirty_bit_2[777] <= 0;lru_counter_1[777] <= 0;lru_counter_2[777] <= 0;tag_1[777] <= 0;tag_2[777] <= 0;cache_mem_1[777] <= 0;cache_mem_2[777] <= 0;
    valid_1[778]  <=   0;valid_2[778]  <=   0;dirty_bit_1[778] <= 0;dirty_bit_2[778] <= 0;lru_counter_1[778] <= 0;lru_counter_2[778] <= 0;tag_1[778] <= 0;tag_2[778] <= 0;cache_mem_1[778] <= 0;cache_mem_2[778] <= 0;
    valid_1[779]  <=   0;valid_2[779]  <=   0;dirty_bit_1[779] <= 0;dirty_bit_2[779] <= 0;lru_counter_1[779] <= 0;lru_counter_2[779] <= 0;tag_1[779] <= 0;tag_2[779] <= 0;cache_mem_1[779] <= 0;cache_mem_2[779] <= 0;
    valid_1[780]  <=   0;valid_2[780]  <=   0;dirty_bit_1[780] <= 0;dirty_bit_2[780] <= 0;lru_counter_1[780] <= 0;lru_counter_2[780] <= 0;tag_1[780] <= 0;tag_2[780] <= 0;cache_mem_1[780] <= 0;cache_mem_2[780] <= 0;
    valid_1[781]  <=   0;valid_2[781]  <=   0;dirty_bit_1[781] <= 0;dirty_bit_2[781] <= 0;lru_counter_1[781] <= 0;lru_counter_2[781] <= 0;tag_1[781] <= 0;tag_2[781] <= 0;cache_mem_1[781] <= 0;cache_mem_2[781] <= 0;
    valid_1[782]  <=   0;valid_2[782]  <=   0;dirty_bit_1[782] <= 0;dirty_bit_2[782] <= 0;lru_counter_1[782] <= 0;lru_counter_2[782] <= 0;tag_1[782] <= 0;tag_2[782] <= 0;cache_mem_1[782] <= 0;cache_mem_2[782] <= 0;
    valid_1[783]  <=   0;valid_2[783]  <=   0;dirty_bit_1[783] <= 0;dirty_bit_2[783] <= 0;lru_counter_1[783] <= 0;lru_counter_2[783] <= 0;tag_1[783] <= 0;tag_2[783] <= 0;cache_mem_1[783] <= 0;cache_mem_2[783] <= 0;
    valid_1[784]  <=   0;valid_2[784]  <=   0;dirty_bit_1[784] <= 0;dirty_bit_2[784] <= 0;lru_counter_1[784] <= 0;lru_counter_2[784] <= 0;tag_1[784] <= 0;tag_2[784] <= 0;cache_mem_1[784] <= 0;cache_mem_2[784] <= 0;
    valid_1[785]  <=   0;valid_2[785]  <=   0;dirty_bit_1[785] <= 0;dirty_bit_2[785] <= 0;lru_counter_1[785] <= 0;lru_counter_2[785] <= 0;tag_1[785] <= 0;tag_2[785] <= 0;cache_mem_1[785] <= 0;cache_mem_2[785] <= 0;
    valid_1[786]  <=   0;valid_2[786]  <=   0;dirty_bit_1[786] <= 0;dirty_bit_2[786] <= 0;lru_counter_1[786] <= 0;lru_counter_2[786] <= 0;tag_1[786] <= 0;tag_2[786] <= 0;cache_mem_1[786] <= 0;cache_mem_2[786] <= 0;
    valid_1[787]  <=   0;valid_2[787]  <=   0;dirty_bit_1[787] <= 0;dirty_bit_2[787] <= 0;lru_counter_1[787] <= 0;lru_counter_2[787] <= 0;tag_1[787] <= 0;tag_2[787] <= 0;cache_mem_1[787] <= 0;cache_mem_2[787] <= 0;
    valid_1[788]  <=   0;valid_2[788]  <=   0;dirty_bit_1[788] <= 0;dirty_bit_2[788] <= 0;lru_counter_1[788] <= 0;lru_counter_2[788] <= 0;tag_1[788] <= 0;tag_2[788] <= 0;cache_mem_1[788] <= 0;cache_mem_2[788] <= 0;
    valid_1[789]  <=   0;valid_2[789]  <=   0;dirty_bit_1[789] <= 0;dirty_bit_2[789] <= 0;lru_counter_1[789] <= 0;lru_counter_2[789] <= 0;tag_1[789] <= 0;tag_2[789] <= 0;cache_mem_1[789] <= 0;cache_mem_2[789] <= 0;
    valid_1[790]  <=   0;valid_2[790]  <=   0;dirty_bit_1[790] <= 0;dirty_bit_2[790] <= 0;lru_counter_1[790] <= 0;lru_counter_2[790] <= 0;tag_1[790] <= 0;tag_2[790] <= 0;cache_mem_1[790] <= 0;cache_mem_2[790] <= 0;
    valid_1[791]  <=   0;valid_2[791]  <=   0;dirty_bit_1[791] <= 0;dirty_bit_2[791] <= 0;lru_counter_1[791] <= 0;lru_counter_2[791] <= 0;tag_1[791] <= 0;tag_2[791] <= 0;cache_mem_1[791] <= 0;cache_mem_2[791] <= 0;
    valid_1[792]  <=   0;valid_2[792]  <=   0;dirty_bit_1[792] <= 0;dirty_bit_2[792] <= 0;lru_counter_1[792] <= 0;lru_counter_2[792] <= 0;tag_1[792] <= 0;tag_2[792] <= 0;cache_mem_1[792] <= 0;cache_mem_2[792] <= 0;
    valid_1[793]  <=   0;valid_2[793]  <=   0;dirty_bit_1[793] <= 0;dirty_bit_2[793] <= 0;lru_counter_1[793] <= 0;lru_counter_2[793] <= 0;tag_1[793] <= 0;tag_2[793] <= 0;cache_mem_1[793] <= 0;cache_mem_2[793] <= 0;
    valid_1[794]  <=   0;valid_2[794]  <=   0;dirty_bit_1[794] <= 0;dirty_bit_2[794] <= 0;lru_counter_1[794] <= 0;lru_counter_2[794] <= 0;tag_1[794] <= 0;tag_2[794] <= 0;cache_mem_1[794] <= 0;cache_mem_2[794] <= 0;
    valid_1[795]  <=   0;valid_2[795]  <=   0;dirty_bit_1[795] <= 0;dirty_bit_2[795] <= 0;lru_counter_1[795] <= 0;lru_counter_2[795] <= 0;tag_1[795] <= 0;tag_2[795] <= 0;cache_mem_1[795] <= 0;cache_mem_2[795] <= 0;
    valid_1[796]  <=   0;valid_2[796]  <=   0;dirty_bit_1[796] <= 0;dirty_bit_2[796] <= 0;lru_counter_1[796] <= 0;lru_counter_2[796] <= 0;tag_1[796] <= 0;tag_2[796] <= 0;cache_mem_1[796] <= 0;cache_mem_2[796] <= 0;
    valid_1[797]  <=   0;valid_2[797]  <=   0;dirty_bit_1[797] <= 0;dirty_bit_2[797] <= 0;lru_counter_1[797] <= 0;lru_counter_2[797] <= 0;tag_1[797] <= 0;tag_2[797] <= 0;cache_mem_1[797] <= 0;cache_mem_2[797] <= 0;
    valid_1[798]  <=   0;valid_2[798]  <=   0;dirty_bit_1[798] <= 0;dirty_bit_2[798] <= 0;lru_counter_1[798] <= 0;lru_counter_2[798] <= 0;tag_1[798] <= 0;tag_2[798] <= 0;cache_mem_1[798] <= 0;cache_mem_2[798] <= 0;
    valid_1[799]  <=   0;valid_2[799]  <=   0;dirty_bit_1[799] <= 0;dirty_bit_2[799] <= 0;lru_counter_1[799] <= 0;lru_counter_2[799] <= 0;tag_1[799] <= 0;tag_2[799] <= 0;cache_mem_1[799] <= 0;cache_mem_2[799] <= 0;
    valid_1[800]  <=   0;valid_2[800]  <=   0;dirty_bit_1[800] <= 0;dirty_bit_2[800] <= 0;lru_counter_1[800] <= 0;lru_counter_2[800] <= 0;tag_1[800] <= 0;tag_2[800] <= 0;cache_mem_1[800] <= 0;cache_mem_2[800] <= 0;
    valid_1[801]  <=   0;valid_2[801]  <=   0;dirty_bit_1[801] <= 0;dirty_bit_2[801] <= 0;lru_counter_1[801] <= 0;lru_counter_2[801] <= 0;tag_1[801] <= 0;tag_2[801] <= 0;cache_mem_1[801] <= 0;cache_mem_2[801] <= 0;
    valid_1[802]  <=   0;valid_2[802]  <=   0;dirty_bit_1[802] <= 0;dirty_bit_2[802] <= 0;lru_counter_1[802] <= 0;lru_counter_2[802] <= 0;tag_1[802] <= 0;tag_2[802] <= 0;cache_mem_1[802] <= 0;cache_mem_2[802] <= 0;
    valid_1[803]  <=   0;valid_2[803]  <=   0;dirty_bit_1[803] <= 0;dirty_bit_2[803] <= 0;lru_counter_1[803] <= 0;lru_counter_2[803] <= 0;tag_1[803] <= 0;tag_2[803] <= 0;cache_mem_1[803] <= 0;cache_mem_2[803] <= 0;
    valid_1[804]  <=   0;valid_2[804]  <=   0;dirty_bit_1[804] <= 0;dirty_bit_2[804] <= 0;lru_counter_1[804] <= 0;lru_counter_2[804] <= 0;tag_1[804] <= 0;tag_2[804] <= 0;cache_mem_1[804] <= 0;cache_mem_2[804] <= 0;
    valid_1[805]  <=   0;valid_2[805]  <=   0;dirty_bit_1[805] <= 0;dirty_bit_2[805] <= 0;lru_counter_1[805] <= 0;lru_counter_2[805] <= 0;tag_1[805] <= 0;tag_2[805] <= 0;cache_mem_1[805] <= 0;cache_mem_2[805] <= 0;
    valid_1[806]  <=   0;valid_2[806]  <=   0;dirty_bit_1[806] <= 0;dirty_bit_2[806] <= 0;lru_counter_1[806] <= 0;lru_counter_2[806] <= 0;tag_1[806] <= 0;tag_2[806] <= 0;cache_mem_1[806] <= 0;cache_mem_2[806] <= 0;
    valid_1[807]  <=   0;valid_2[807]  <=   0;dirty_bit_1[807] <= 0;dirty_bit_2[807] <= 0;lru_counter_1[807] <= 0;lru_counter_2[807] <= 0;tag_1[807] <= 0;tag_2[807] <= 0;cache_mem_1[807] <= 0;cache_mem_2[807] <= 0;
    valid_1[808]  <=   0;valid_2[808]  <=   0;dirty_bit_1[808] <= 0;dirty_bit_2[808] <= 0;lru_counter_1[808] <= 0;lru_counter_2[808] <= 0;tag_1[808] <= 0;tag_2[808] <= 0;cache_mem_1[808] <= 0;cache_mem_2[808] <= 0;
    valid_1[809]  <=   0;valid_2[809]  <=   0;dirty_bit_1[809] <= 0;dirty_bit_2[809] <= 0;lru_counter_1[809] <= 0;lru_counter_2[809] <= 0;tag_1[809] <= 0;tag_2[809] <= 0;cache_mem_1[809] <= 0;cache_mem_2[809] <= 0;
    valid_1[810]  <=   0;valid_2[810]  <=   0;dirty_bit_1[810] <= 0;dirty_bit_2[810] <= 0;lru_counter_1[810] <= 0;lru_counter_2[810] <= 0;tag_1[810] <= 0;tag_2[810] <= 0;cache_mem_1[810] <= 0;cache_mem_2[810] <= 0;
    valid_1[811]  <=   0;valid_2[811]  <=   0;dirty_bit_1[811] <= 0;dirty_bit_2[811] <= 0;lru_counter_1[811] <= 0;lru_counter_2[811] <= 0;tag_1[811] <= 0;tag_2[811] <= 0;cache_mem_1[811] <= 0;cache_mem_2[811] <= 0;
    valid_1[812]  <=   0;valid_2[812]  <=   0;dirty_bit_1[812] <= 0;dirty_bit_2[812] <= 0;lru_counter_1[812] <= 0;lru_counter_2[812] <= 0;tag_1[812] <= 0;tag_2[812] <= 0;cache_mem_1[812] <= 0;cache_mem_2[812] <= 0;
    valid_1[813]  <=   0;valid_2[813]  <=   0;dirty_bit_1[813] <= 0;dirty_bit_2[813] <= 0;lru_counter_1[813] <= 0;lru_counter_2[813] <= 0;tag_1[813] <= 0;tag_2[813] <= 0;cache_mem_1[813] <= 0;cache_mem_2[813] <= 0;
    valid_1[814]  <=   0;valid_2[814]  <=   0;dirty_bit_1[814] <= 0;dirty_bit_2[814] <= 0;lru_counter_1[814] <= 0;lru_counter_2[814] <= 0;tag_1[814] <= 0;tag_2[814] <= 0;cache_mem_1[814] <= 0;cache_mem_2[814] <= 0;
    valid_1[815]  <=   0;valid_2[815]  <=   0;dirty_bit_1[815] <= 0;dirty_bit_2[815] <= 0;lru_counter_1[815] <= 0;lru_counter_2[815] <= 0;tag_1[815] <= 0;tag_2[815] <= 0;cache_mem_1[815] <= 0;cache_mem_2[815] <= 0;
    valid_1[816]  <=   0;valid_2[816]  <=   0;dirty_bit_1[816] <= 0;dirty_bit_2[816] <= 0;lru_counter_1[816] <= 0;lru_counter_2[816] <= 0;tag_1[816] <= 0;tag_2[816] <= 0;cache_mem_1[816] <= 0;cache_mem_2[816] <= 0;
    valid_1[817]  <=   0;valid_2[817]  <=   0;dirty_bit_1[817] <= 0;dirty_bit_2[817] <= 0;lru_counter_1[817] <= 0;lru_counter_2[817] <= 0;tag_1[817] <= 0;tag_2[817] <= 0;cache_mem_1[817] <= 0;cache_mem_2[817] <= 0;
    valid_1[818]  <=   0;valid_2[818]  <=   0;dirty_bit_1[818] <= 0;dirty_bit_2[818] <= 0;lru_counter_1[818] <= 0;lru_counter_2[818] <= 0;tag_1[818] <= 0;tag_2[818] <= 0;cache_mem_1[818] <= 0;cache_mem_2[818] <= 0;
    valid_1[819]  <=   0;valid_2[819]  <=   0;dirty_bit_1[819] <= 0;dirty_bit_2[819] <= 0;lru_counter_1[819] <= 0;lru_counter_2[819] <= 0;tag_1[819] <= 0;tag_2[819] <= 0;cache_mem_1[819] <= 0;cache_mem_2[819] <= 0;
    valid_1[820]  <=   0;valid_2[820]  <=   0;dirty_bit_1[820] <= 0;dirty_bit_2[820] <= 0;lru_counter_1[820] <= 0;lru_counter_2[820] <= 0;tag_1[820] <= 0;tag_2[820] <= 0;cache_mem_1[820] <= 0;cache_mem_2[820] <= 0;
    valid_1[821]  <=   0;valid_2[821]  <=   0;dirty_bit_1[821] <= 0;dirty_bit_2[821] <= 0;lru_counter_1[821] <= 0;lru_counter_2[821] <= 0;tag_1[821] <= 0;tag_2[821] <= 0;cache_mem_1[821] <= 0;cache_mem_2[821] <= 0;
    valid_1[822]  <=   0;valid_2[822]  <=   0;dirty_bit_1[822] <= 0;dirty_bit_2[822] <= 0;lru_counter_1[822] <= 0;lru_counter_2[822] <= 0;tag_1[822] <= 0;tag_2[822] <= 0;cache_mem_1[822] <= 0;cache_mem_2[822] <= 0;
    valid_1[823]  <=   0;valid_2[823]  <=   0;dirty_bit_1[823] <= 0;dirty_bit_2[823] <= 0;lru_counter_1[823] <= 0;lru_counter_2[823] <= 0;tag_1[823] <= 0;tag_2[823] <= 0;cache_mem_1[823] <= 0;cache_mem_2[823] <= 0;
    valid_1[824]  <=   0;valid_2[824]  <=   0;dirty_bit_1[824] <= 0;dirty_bit_2[824] <= 0;lru_counter_1[824] <= 0;lru_counter_2[824] <= 0;tag_1[824] <= 0;tag_2[824] <= 0;cache_mem_1[824] <= 0;cache_mem_2[824] <= 0;
    valid_1[825]  <=   0;valid_2[825]  <=   0;dirty_bit_1[825] <= 0;dirty_bit_2[825] <= 0;lru_counter_1[825] <= 0;lru_counter_2[825] <= 0;tag_1[825] <= 0;tag_2[825] <= 0;cache_mem_1[825] <= 0;cache_mem_2[825] <= 0;
    valid_1[826]  <=   0;valid_2[826]  <=   0;dirty_bit_1[826] <= 0;dirty_bit_2[826] <= 0;lru_counter_1[826] <= 0;lru_counter_2[826] <= 0;tag_1[826] <= 0;tag_2[826] <= 0;cache_mem_1[826] <= 0;cache_mem_2[826] <= 0;
    valid_1[827]  <=   0;valid_2[827]  <=   0;dirty_bit_1[827] <= 0;dirty_bit_2[827] <= 0;lru_counter_1[827] <= 0;lru_counter_2[827] <= 0;tag_1[827] <= 0;tag_2[827] <= 0;cache_mem_1[827] <= 0;cache_mem_2[827] <= 0;
    valid_1[828]  <=   0;valid_2[828]  <=   0;dirty_bit_1[828] <= 0;dirty_bit_2[828] <= 0;lru_counter_1[828] <= 0;lru_counter_2[828] <= 0;tag_1[828] <= 0;tag_2[828] <= 0;cache_mem_1[828] <= 0;cache_mem_2[828] <= 0;
    valid_1[829]  <=   0;valid_2[829]  <=   0;dirty_bit_1[829] <= 0;dirty_bit_2[829] <= 0;lru_counter_1[829] <= 0;lru_counter_2[829] <= 0;tag_1[829] <= 0;tag_2[829] <= 0;cache_mem_1[829] <= 0;cache_mem_2[829] <= 0;
    valid_1[830]  <=   0;valid_2[830]  <=   0;dirty_bit_1[830] <= 0;dirty_bit_2[830] <= 0;lru_counter_1[830] <= 0;lru_counter_2[830] <= 0;tag_1[830] <= 0;tag_2[830] <= 0;cache_mem_1[830] <= 0;cache_mem_2[830] <= 0;
    valid_1[831]  <=   0;valid_2[831]  <=   0;dirty_bit_1[831] <= 0;dirty_bit_2[831] <= 0;lru_counter_1[831] <= 0;lru_counter_2[831] <= 0;tag_1[831] <= 0;tag_2[831] <= 0;cache_mem_1[831] <= 0;cache_mem_2[831] <= 0;
    valid_1[832]  <=   0;valid_2[832]  <=   0;dirty_bit_1[832] <= 0;dirty_bit_2[832] <= 0;lru_counter_1[832] <= 0;lru_counter_2[832] <= 0;tag_1[832] <= 0;tag_2[832] <= 0;cache_mem_1[832] <= 0;cache_mem_2[832] <= 0;
    valid_1[833]  <=   0;valid_2[833]  <=   0;dirty_bit_1[833] <= 0;dirty_bit_2[833] <= 0;lru_counter_1[833] <= 0;lru_counter_2[833] <= 0;tag_1[833] <= 0;tag_2[833] <= 0;cache_mem_1[833] <= 0;cache_mem_2[833] <= 0;
    valid_1[834]  <=   0;valid_2[834]  <=   0;dirty_bit_1[834] <= 0;dirty_bit_2[834] <= 0;lru_counter_1[834] <= 0;lru_counter_2[834] <= 0;tag_1[834] <= 0;tag_2[834] <= 0;cache_mem_1[834] <= 0;cache_mem_2[834] <= 0;
    valid_1[835]  <=   0;valid_2[835]  <=   0;dirty_bit_1[835] <= 0;dirty_bit_2[835] <= 0;lru_counter_1[835] <= 0;lru_counter_2[835] <= 0;tag_1[835] <= 0;tag_2[835] <= 0;cache_mem_1[835] <= 0;cache_mem_2[835] <= 0;
    valid_1[836]  <=   0;valid_2[836]  <=   0;dirty_bit_1[836] <= 0;dirty_bit_2[836] <= 0;lru_counter_1[836] <= 0;lru_counter_2[836] <= 0;tag_1[836] <= 0;tag_2[836] <= 0;cache_mem_1[836] <= 0;cache_mem_2[836] <= 0;
    valid_1[837]  <=   0;valid_2[837]  <=   0;dirty_bit_1[837] <= 0;dirty_bit_2[837] <= 0;lru_counter_1[837] <= 0;lru_counter_2[837] <= 0;tag_1[837] <= 0;tag_2[837] <= 0;cache_mem_1[837] <= 0;cache_mem_2[837] <= 0;
    valid_1[838]  <=   0;valid_2[838]  <=   0;dirty_bit_1[838] <= 0;dirty_bit_2[838] <= 0;lru_counter_1[838] <= 0;lru_counter_2[838] <= 0;tag_1[838] <= 0;tag_2[838] <= 0;cache_mem_1[838] <= 0;cache_mem_2[838] <= 0;
    valid_1[839]  <=   0;valid_2[839]  <=   0;dirty_bit_1[839] <= 0;dirty_bit_2[839] <= 0;lru_counter_1[839] <= 0;lru_counter_2[839] <= 0;tag_1[839] <= 0;tag_2[839] <= 0;cache_mem_1[839] <= 0;cache_mem_2[839] <= 0;
    valid_1[840]  <=   0;valid_2[840]  <=   0;dirty_bit_1[840] <= 0;dirty_bit_2[840] <= 0;lru_counter_1[840] <= 0;lru_counter_2[840] <= 0;tag_1[840] <= 0;tag_2[840] <= 0;cache_mem_1[840] <= 0;cache_mem_2[840] <= 0;
    valid_1[841]  <=   0;valid_2[841]  <=   0;dirty_bit_1[841] <= 0;dirty_bit_2[841] <= 0;lru_counter_1[841] <= 0;lru_counter_2[841] <= 0;tag_1[841] <= 0;tag_2[841] <= 0;cache_mem_1[841] <= 0;cache_mem_2[841] <= 0;
    valid_1[842]  <=   0;valid_2[842]  <=   0;dirty_bit_1[842] <= 0;dirty_bit_2[842] <= 0;lru_counter_1[842] <= 0;lru_counter_2[842] <= 0;tag_1[842] <= 0;tag_2[842] <= 0;cache_mem_1[842] <= 0;cache_mem_2[842] <= 0;
    valid_1[843]  <=   0;valid_2[843]  <=   0;dirty_bit_1[843] <= 0;dirty_bit_2[843] <= 0;lru_counter_1[843] <= 0;lru_counter_2[843] <= 0;tag_1[843] <= 0;tag_2[843] <= 0;cache_mem_1[843] <= 0;cache_mem_2[843] <= 0;
    valid_1[844]  <=   0;valid_2[844]  <=   0;dirty_bit_1[844] <= 0;dirty_bit_2[844] <= 0;lru_counter_1[844] <= 0;lru_counter_2[844] <= 0;tag_1[844] <= 0;tag_2[844] <= 0;cache_mem_1[844] <= 0;cache_mem_2[844] <= 0;
    valid_1[845]  <=   0;valid_2[845]  <=   0;dirty_bit_1[845] <= 0;dirty_bit_2[845] <= 0;lru_counter_1[845] <= 0;lru_counter_2[845] <= 0;tag_1[845] <= 0;tag_2[845] <= 0;cache_mem_1[845] <= 0;cache_mem_2[845] <= 0;
    valid_1[846]  <=   0;valid_2[846]  <=   0;dirty_bit_1[846] <= 0;dirty_bit_2[846] <= 0;lru_counter_1[846] <= 0;lru_counter_2[846] <= 0;tag_1[846] <= 0;tag_2[846] <= 0;cache_mem_1[846] <= 0;cache_mem_2[846] <= 0;
    valid_1[847]  <=   0;valid_2[847]  <=   0;dirty_bit_1[847] <= 0;dirty_bit_2[847] <= 0;lru_counter_1[847] <= 0;lru_counter_2[847] <= 0;tag_1[847] <= 0;tag_2[847] <= 0;cache_mem_1[847] <= 0;cache_mem_2[847] <= 0;
    valid_1[848]  <=   0;valid_2[848]  <=   0;dirty_bit_1[848] <= 0;dirty_bit_2[848] <= 0;lru_counter_1[848] <= 0;lru_counter_2[848] <= 0;tag_1[848] <= 0;tag_2[848] <= 0;cache_mem_1[848] <= 0;cache_mem_2[848] <= 0;
    valid_1[849]  <=   0;valid_2[849]  <=   0;dirty_bit_1[849] <= 0;dirty_bit_2[849] <= 0;lru_counter_1[849] <= 0;lru_counter_2[849] <= 0;tag_1[849] <= 0;tag_2[849] <= 0;cache_mem_1[849] <= 0;cache_mem_2[849] <= 0;
    valid_1[850]  <=   0;valid_2[850]  <=   0;dirty_bit_1[850] <= 0;dirty_bit_2[850] <= 0;lru_counter_1[850] <= 0;lru_counter_2[850] <= 0;tag_1[850] <= 0;tag_2[850] <= 0;cache_mem_1[850] <= 0;cache_mem_2[850] <= 0;
    valid_1[851]  <=   0;valid_2[851]  <=   0;dirty_bit_1[851] <= 0;dirty_bit_2[851] <= 0;lru_counter_1[851] <= 0;lru_counter_2[851] <= 0;tag_1[851] <= 0;tag_2[851] <= 0;cache_mem_1[851] <= 0;cache_mem_2[851] <= 0;
    valid_1[852]  <=   0;valid_2[852]  <=   0;dirty_bit_1[852] <= 0;dirty_bit_2[852] <= 0;lru_counter_1[852] <= 0;lru_counter_2[852] <= 0;tag_1[852] <= 0;tag_2[852] <= 0;cache_mem_1[852] <= 0;cache_mem_2[852] <= 0;
    valid_1[853]  <=   0;valid_2[853]  <=   0;dirty_bit_1[853] <= 0;dirty_bit_2[853] <= 0;lru_counter_1[853] <= 0;lru_counter_2[853] <= 0;tag_1[853] <= 0;tag_2[853] <= 0;cache_mem_1[853] <= 0;cache_mem_2[853] <= 0;
    valid_1[854]  <=   0;valid_2[854]  <=   0;dirty_bit_1[854] <= 0;dirty_bit_2[854] <= 0;lru_counter_1[854] <= 0;lru_counter_2[854] <= 0;tag_1[854] <= 0;tag_2[854] <= 0;cache_mem_1[854] <= 0;cache_mem_2[854] <= 0;
    valid_1[855]  <=   0;valid_2[855]  <=   0;dirty_bit_1[855] <= 0;dirty_bit_2[855] <= 0;lru_counter_1[855] <= 0;lru_counter_2[855] <= 0;tag_1[855] <= 0;tag_2[855] <= 0;cache_mem_1[855] <= 0;cache_mem_2[855] <= 0;
    valid_1[856]  <=   0;valid_2[856]  <=   0;dirty_bit_1[856] <= 0;dirty_bit_2[856] <= 0;lru_counter_1[856] <= 0;lru_counter_2[856] <= 0;tag_1[856] <= 0;tag_2[856] <= 0;cache_mem_1[856] <= 0;cache_mem_2[856] <= 0;
    valid_1[857]  <=   0;valid_2[857]  <=   0;dirty_bit_1[857] <= 0;dirty_bit_2[857] <= 0;lru_counter_1[857] <= 0;lru_counter_2[857] <= 0;tag_1[857] <= 0;tag_2[857] <= 0;cache_mem_1[857] <= 0;cache_mem_2[857] <= 0;
    valid_1[858]  <=   0;valid_2[858]  <=   0;dirty_bit_1[858] <= 0;dirty_bit_2[858] <= 0;lru_counter_1[858] <= 0;lru_counter_2[858] <= 0;tag_1[858] <= 0;tag_2[858] <= 0;cache_mem_1[858] <= 0;cache_mem_2[858] <= 0;
    valid_1[859]  <=   0;valid_2[859]  <=   0;dirty_bit_1[859] <= 0;dirty_bit_2[859] <= 0;lru_counter_1[859] <= 0;lru_counter_2[859] <= 0;tag_1[859] <= 0;tag_2[859] <= 0;cache_mem_1[859] <= 0;cache_mem_2[859] <= 0;
    valid_1[860]  <=   0;valid_2[860]  <=   0;dirty_bit_1[860] <= 0;dirty_bit_2[860] <= 0;lru_counter_1[860] <= 0;lru_counter_2[860] <= 0;tag_1[860] <= 0;tag_2[860] <= 0;cache_mem_1[860] <= 0;cache_mem_2[860] <= 0;
    valid_1[861]  <=   0;valid_2[861]  <=   0;dirty_bit_1[861] <= 0;dirty_bit_2[861] <= 0;lru_counter_1[861] <= 0;lru_counter_2[861] <= 0;tag_1[861] <= 0;tag_2[861] <= 0;cache_mem_1[861] <= 0;cache_mem_2[861] <= 0;
    valid_1[862]  <=   0;valid_2[862]  <=   0;dirty_bit_1[862] <= 0;dirty_bit_2[862] <= 0;lru_counter_1[862] <= 0;lru_counter_2[862] <= 0;tag_1[862] <= 0;tag_2[862] <= 0;cache_mem_1[862] <= 0;cache_mem_2[862] <= 0;
    valid_1[863]  <=   0;valid_2[863]  <=   0;dirty_bit_1[863] <= 0;dirty_bit_2[863] <= 0;lru_counter_1[863] <= 0;lru_counter_2[863] <= 0;tag_1[863] <= 0;tag_2[863] <= 0;cache_mem_1[863] <= 0;cache_mem_2[863] <= 0;
    valid_1[864]  <=   0;valid_2[864]  <=   0;dirty_bit_1[864] <= 0;dirty_bit_2[864] <= 0;lru_counter_1[864] <= 0;lru_counter_2[864] <= 0;tag_1[864] <= 0;tag_2[864] <= 0;cache_mem_1[864] <= 0;cache_mem_2[864] <= 0;
    valid_1[865]  <=   0;valid_2[865]  <=   0;dirty_bit_1[865] <= 0;dirty_bit_2[865] <= 0;lru_counter_1[865] <= 0;lru_counter_2[865] <= 0;tag_1[865] <= 0;tag_2[865] <= 0;cache_mem_1[865] <= 0;cache_mem_2[865] <= 0;
    valid_1[866]  <=   0;valid_2[866]  <=   0;dirty_bit_1[866] <= 0;dirty_bit_2[866] <= 0;lru_counter_1[866] <= 0;lru_counter_2[866] <= 0;tag_1[866] <= 0;tag_2[866] <= 0;cache_mem_1[866] <= 0;cache_mem_2[866] <= 0;
    valid_1[867]  <=   0;valid_2[867]  <=   0;dirty_bit_1[867] <= 0;dirty_bit_2[867] <= 0;lru_counter_1[867] <= 0;lru_counter_2[867] <= 0;tag_1[867] <= 0;tag_2[867] <= 0;cache_mem_1[867] <= 0;cache_mem_2[867] <= 0;
    valid_1[868]  <=   0;valid_2[868]  <=   0;dirty_bit_1[868] <= 0;dirty_bit_2[868] <= 0;lru_counter_1[868] <= 0;lru_counter_2[868] <= 0;tag_1[868] <= 0;tag_2[868] <= 0;cache_mem_1[868] <= 0;cache_mem_2[868] <= 0;
    valid_1[869]  <=   0;valid_2[869]  <=   0;dirty_bit_1[869] <= 0;dirty_bit_2[869] <= 0;lru_counter_1[869] <= 0;lru_counter_2[869] <= 0;tag_1[869] <= 0;tag_2[869] <= 0;cache_mem_1[869] <= 0;cache_mem_2[869] <= 0;
    valid_1[870]  <=   0;valid_2[870]  <=   0;dirty_bit_1[870] <= 0;dirty_bit_2[870] <= 0;lru_counter_1[870] <= 0;lru_counter_2[870] <= 0;tag_1[870] <= 0;tag_2[870] <= 0;cache_mem_1[870] <= 0;cache_mem_2[870] <= 0;
    valid_1[871]  <=   0;valid_2[871]  <=   0;dirty_bit_1[871] <= 0;dirty_bit_2[871] <= 0;lru_counter_1[871] <= 0;lru_counter_2[871] <= 0;tag_1[871] <= 0;tag_2[871] <= 0;cache_mem_1[871] <= 0;cache_mem_2[871] <= 0;
    valid_1[872]  <=   0;valid_2[872]  <=   0;dirty_bit_1[872] <= 0;dirty_bit_2[872] <= 0;lru_counter_1[872] <= 0;lru_counter_2[872] <= 0;tag_1[872] <= 0;tag_2[872] <= 0;cache_mem_1[872] <= 0;cache_mem_2[872] <= 0;
    valid_1[873]  <=   0;valid_2[873]  <=   0;dirty_bit_1[873] <= 0;dirty_bit_2[873] <= 0;lru_counter_1[873] <= 0;lru_counter_2[873] <= 0;tag_1[873] <= 0;tag_2[873] <= 0;cache_mem_1[873] <= 0;cache_mem_2[873] <= 0;
    valid_1[874]  <=   0;valid_2[874]  <=   0;dirty_bit_1[874] <= 0;dirty_bit_2[874] <= 0;lru_counter_1[874] <= 0;lru_counter_2[874] <= 0;tag_1[874] <= 0;tag_2[874] <= 0;cache_mem_1[874] <= 0;cache_mem_2[874] <= 0;
    valid_1[875]  <=   0;valid_2[875]  <=   0;dirty_bit_1[875] <= 0;dirty_bit_2[875] <= 0;lru_counter_1[875] <= 0;lru_counter_2[875] <= 0;tag_1[875] <= 0;tag_2[875] <= 0;cache_mem_1[875] <= 0;cache_mem_2[875] <= 0;
    valid_1[876]  <=   0;valid_2[876]  <=   0;dirty_bit_1[876] <= 0;dirty_bit_2[876] <= 0;lru_counter_1[876] <= 0;lru_counter_2[876] <= 0;tag_1[876] <= 0;tag_2[876] <= 0;cache_mem_1[876] <= 0;cache_mem_2[876] <= 0;
    valid_1[877]  <=   0;valid_2[877]  <=   0;dirty_bit_1[877] <= 0;dirty_bit_2[877] <= 0;lru_counter_1[877] <= 0;lru_counter_2[877] <= 0;tag_1[877] <= 0;tag_2[877] <= 0;cache_mem_1[877] <= 0;cache_mem_2[877] <= 0;
    valid_1[878]  <=   0;valid_2[878]  <=   0;dirty_bit_1[878] <= 0;dirty_bit_2[878] <= 0;lru_counter_1[878] <= 0;lru_counter_2[878] <= 0;tag_1[878] <= 0;tag_2[878] <= 0;cache_mem_1[878] <= 0;cache_mem_2[878] <= 0;
    valid_1[879]  <=   0;valid_2[879]  <=   0;dirty_bit_1[879] <= 0;dirty_bit_2[879] <= 0;lru_counter_1[879] <= 0;lru_counter_2[879] <= 0;tag_1[879] <= 0;tag_2[879] <= 0;cache_mem_1[879] <= 0;cache_mem_2[879] <= 0;
    valid_1[880]  <=   0;valid_2[880]  <=   0;dirty_bit_1[880] <= 0;dirty_bit_2[880] <= 0;lru_counter_1[880] <= 0;lru_counter_2[880] <= 0;tag_1[880] <= 0;tag_2[880] <= 0;cache_mem_1[880] <= 0;cache_mem_2[880] <= 0;
    valid_1[881]  <=   0;valid_2[881]  <=   0;dirty_bit_1[881] <= 0;dirty_bit_2[881] <= 0;lru_counter_1[881] <= 0;lru_counter_2[881] <= 0;tag_1[881] <= 0;tag_2[881] <= 0;cache_mem_1[881] <= 0;cache_mem_2[881] <= 0;
    valid_1[882]  <=   0;valid_2[882]  <=   0;dirty_bit_1[882] <= 0;dirty_bit_2[882] <= 0;lru_counter_1[882] <= 0;lru_counter_2[882] <= 0;tag_1[882] <= 0;tag_2[882] <= 0;cache_mem_1[882] <= 0;cache_mem_2[882] <= 0;
    valid_1[883]  <=   0;valid_2[883]  <=   0;dirty_bit_1[883] <= 0;dirty_bit_2[883] <= 0;lru_counter_1[883] <= 0;lru_counter_2[883] <= 0;tag_1[883] <= 0;tag_2[883] <= 0;cache_mem_1[883] <= 0;cache_mem_2[883] <= 0;
    valid_1[884]  <=   0;valid_2[884]  <=   0;dirty_bit_1[884] <= 0;dirty_bit_2[884] <= 0;lru_counter_1[884] <= 0;lru_counter_2[884] <= 0;tag_1[884] <= 0;tag_2[884] <= 0;cache_mem_1[884] <= 0;cache_mem_2[884] <= 0;
    valid_1[885]  <=   0;valid_2[885]  <=   0;dirty_bit_1[885] <= 0;dirty_bit_2[885] <= 0;lru_counter_1[885] <= 0;lru_counter_2[885] <= 0;tag_1[885] <= 0;tag_2[885] <= 0;cache_mem_1[885] <= 0;cache_mem_2[885] <= 0;
    valid_1[886]  <=   0;valid_2[886]  <=   0;dirty_bit_1[886] <= 0;dirty_bit_2[886] <= 0;lru_counter_1[886] <= 0;lru_counter_2[886] <= 0;tag_1[886] <= 0;tag_2[886] <= 0;cache_mem_1[886] <= 0;cache_mem_2[886] <= 0;
    valid_1[887]  <=   0;valid_2[887]  <=   0;dirty_bit_1[887] <= 0;dirty_bit_2[887] <= 0;lru_counter_1[887] <= 0;lru_counter_2[887] <= 0;tag_1[887] <= 0;tag_2[887] <= 0;cache_mem_1[887] <= 0;cache_mem_2[887] <= 0;
    valid_1[888]  <=   0;valid_2[888]  <=   0;dirty_bit_1[888] <= 0;dirty_bit_2[888] <= 0;lru_counter_1[888] <= 0;lru_counter_2[888] <= 0;tag_1[888] <= 0;tag_2[888] <= 0;cache_mem_1[888] <= 0;cache_mem_2[888] <= 0;
    valid_1[889]  <=   0;valid_2[889]  <=   0;dirty_bit_1[889] <= 0;dirty_bit_2[889] <= 0;lru_counter_1[889] <= 0;lru_counter_2[889] <= 0;tag_1[889] <= 0;tag_2[889] <= 0;cache_mem_1[889] <= 0;cache_mem_2[889] <= 0;
    valid_1[890]  <=   0;valid_2[890]  <=   0;dirty_bit_1[890] <= 0;dirty_bit_2[890] <= 0;lru_counter_1[890] <= 0;lru_counter_2[890] <= 0;tag_1[890] <= 0;tag_2[890] <= 0;cache_mem_1[890] <= 0;cache_mem_2[890] <= 0;
    valid_1[891]  <=   0;valid_2[891]  <=   0;dirty_bit_1[891] <= 0;dirty_bit_2[891] <= 0;lru_counter_1[891] <= 0;lru_counter_2[891] <= 0;tag_1[891] <= 0;tag_2[891] <= 0;cache_mem_1[891] <= 0;cache_mem_2[891] <= 0;
    valid_1[892]  <=   0;valid_2[892]  <=   0;dirty_bit_1[892] <= 0;dirty_bit_2[892] <= 0;lru_counter_1[892] <= 0;lru_counter_2[892] <= 0;tag_1[892] <= 0;tag_2[892] <= 0;cache_mem_1[892] <= 0;cache_mem_2[892] <= 0;
    valid_1[893]  <=   0;valid_2[893]  <=   0;dirty_bit_1[893] <= 0;dirty_bit_2[893] <= 0;lru_counter_1[893] <= 0;lru_counter_2[893] <= 0;tag_1[893] <= 0;tag_2[893] <= 0;cache_mem_1[893] <= 0;cache_mem_2[893] <= 0;
    valid_1[894]  <=   0;valid_2[894]  <=   0;dirty_bit_1[894] <= 0;dirty_bit_2[894] <= 0;lru_counter_1[894] <= 0;lru_counter_2[894] <= 0;tag_1[894] <= 0;tag_2[894] <= 0;cache_mem_1[894] <= 0;cache_mem_2[894] <= 0;
    valid_1[895]  <=   0;valid_2[895]  <=   0;dirty_bit_1[895] <= 0;dirty_bit_2[895] <= 0;lru_counter_1[895] <= 0;lru_counter_2[895] <= 0;tag_1[895] <= 0;tag_2[895] <= 0;cache_mem_1[895] <= 0;cache_mem_2[895] <= 0;
    valid_1[896]  <=   0;valid_2[896]  <=   0;dirty_bit_1[896] <= 0;dirty_bit_2[896] <= 0;lru_counter_1[896] <= 0;lru_counter_2[896] <= 0;tag_1[896] <= 0;tag_2[896] <= 0;cache_mem_1[896] <= 0;cache_mem_2[896] <= 0;
    valid_1[897]  <=   0;valid_2[897]  <=   0;dirty_bit_1[897] <= 0;dirty_bit_2[897] <= 0;lru_counter_1[897] <= 0;lru_counter_2[897] <= 0;tag_1[897] <= 0;tag_2[897] <= 0;cache_mem_1[897] <= 0;cache_mem_2[897] <= 0;
    valid_1[898]  <=   0;valid_2[898]  <=   0;dirty_bit_1[898] <= 0;dirty_bit_2[898] <= 0;lru_counter_1[898] <= 0;lru_counter_2[898] <= 0;tag_1[898] <= 0;tag_2[898] <= 0;cache_mem_1[898] <= 0;cache_mem_2[898] <= 0;
    valid_1[899]  <=   0;valid_2[899]  <=   0;dirty_bit_1[899] <= 0;dirty_bit_2[899] <= 0;lru_counter_1[899] <= 0;lru_counter_2[899] <= 0;tag_1[899] <= 0;tag_2[899] <= 0;cache_mem_1[899] <= 0;cache_mem_2[899] <= 0;
    valid_1[900]  <=   0;valid_2[900]  <=   0;dirty_bit_1[900] <= 0;dirty_bit_2[900] <= 0;lru_counter_1[900] <= 0;lru_counter_2[900] <= 0;tag_1[900] <= 0;tag_2[900] <= 0;cache_mem_1[900] <= 0;cache_mem_2[900] <= 0;
    valid_1[901]  <=   0;valid_2[901]  <=   0;dirty_bit_1[901] <= 0;dirty_bit_2[901] <= 0;lru_counter_1[901] <= 0;lru_counter_2[901] <= 0;tag_1[901] <= 0;tag_2[901] <= 0;cache_mem_1[901] <= 0;cache_mem_2[901] <= 0;
    valid_1[902]  <=   0;valid_2[902]  <=   0;dirty_bit_1[902] <= 0;dirty_bit_2[902] <= 0;lru_counter_1[902] <= 0;lru_counter_2[902] <= 0;tag_1[902] <= 0;tag_2[902] <= 0;cache_mem_1[902] <= 0;cache_mem_2[902] <= 0;
    valid_1[903]  <=   0;valid_2[903]  <=   0;dirty_bit_1[903] <= 0;dirty_bit_2[903] <= 0;lru_counter_1[903] <= 0;lru_counter_2[903] <= 0;tag_1[903] <= 0;tag_2[903] <= 0;cache_mem_1[903] <= 0;cache_mem_2[903] <= 0;
    valid_1[904]  <=   0;valid_2[904]  <=   0;dirty_bit_1[904] <= 0;dirty_bit_2[904] <= 0;lru_counter_1[904] <= 0;lru_counter_2[904] <= 0;tag_1[904] <= 0;tag_2[904] <= 0;cache_mem_1[904] <= 0;cache_mem_2[904] <= 0;
    valid_1[905]  <=   0;valid_2[905]  <=   0;dirty_bit_1[905] <= 0;dirty_bit_2[905] <= 0;lru_counter_1[905] <= 0;lru_counter_2[905] <= 0;tag_1[905] <= 0;tag_2[905] <= 0;cache_mem_1[905] <= 0;cache_mem_2[905] <= 0;
    valid_1[906]  <=   0;valid_2[906]  <=   0;dirty_bit_1[906] <= 0;dirty_bit_2[906] <= 0;lru_counter_1[906] <= 0;lru_counter_2[906] <= 0;tag_1[906] <= 0;tag_2[906] <= 0;cache_mem_1[906] <= 0;cache_mem_2[906] <= 0;
    valid_1[907]  <=   0;valid_2[907]  <=   0;dirty_bit_1[907] <= 0;dirty_bit_2[907] <= 0;lru_counter_1[907] <= 0;lru_counter_2[907] <= 0;tag_1[907] <= 0;tag_2[907] <= 0;cache_mem_1[907] <= 0;cache_mem_2[907] <= 0;
    valid_1[908]  <=   0;valid_2[908]  <=   0;dirty_bit_1[908] <= 0;dirty_bit_2[908] <= 0;lru_counter_1[908] <= 0;lru_counter_2[908] <= 0;tag_1[908] <= 0;tag_2[908] <= 0;cache_mem_1[908] <= 0;cache_mem_2[908] <= 0;
    valid_1[909]  <=   0;valid_2[909]  <=   0;dirty_bit_1[909] <= 0;dirty_bit_2[909] <= 0;lru_counter_1[909] <= 0;lru_counter_2[909] <= 0;tag_1[909] <= 0;tag_2[909] <= 0;cache_mem_1[909] <= 0;cache_mem_2[909] <= 0;
    valid_1[910]  <=   0;valid_2[910]  <=   0;dirty_bit_1[910] <= 0;dirty_bit_2[910] <= 0;lru_counter_1[910] <= 0;lru_counter_2[910] <= 0;tag_1[910] <= 0;tag_2[910] <= 0;cache_mem_1[910] <= 0;cache_mem_2[910] <= 0;
    valid_1[911]  <=   0;valid_2[911]  <=   0;dirty_bit_1[911] <= 0;dirty_bit_2[911] <= 0;lru_counter_1[911] <= 0;lru_counter_2[911] <= 0;tag_1[911] <= 0;tag_2[911] <= 0;cache_mem_1[911] <= 0;cache_mem_2[911] <= 0;
    valid_1[912]  <=   0;valid_2[912]  <=   0;dirty_bit_1[912] <= 0;dirty_bit_2[912] <= 0;lru_counter_1[912] <= 0;lru_counter_2[912] <= 0;tag_1[912] <= 0;tag_2[912] <= 0;cache_mem_1[912] <= 0;cache_mem_2[912] <= 0;
    valid_1[913]  <=   0;valid_2[913]  <=   0;dirty_bit_1[913] <= 0;dirty_bit_2[913] <= 0;lru_counter_1[913] <= 0;lru_counter_2[913] <= 0;tag_1[913] <= 0;tag_2[913] <= 0;cache_mem_1[913] <= 0;cache_mem_2[913] <= 0;
    valid_1[914]  <=   0;valid_2[914]  <=   0;dirty_bit_1[914] <= 0;dirty_bit_2[914] <= 0;lru_counter_1[914] <= 0;lru_counter_2[914] <= 0;tag_1[914] <= 0;tag_2[914] <= 0;cache_mem_1[914] <= 0;cache_mem_2[914] <= 0;
    valid_1[915]  <=   0;valid_2[915]  <=   0;dirty_bit_1[915] <= 0;dirty_bit_2[915] <= 0;lru_counter_1[915] <= 0;lru_counter_2[915] <= 0;tag_1[915] <= 0;tag_2[915] <= 0;cache_mem_1[915] <= 0;cache_mem_2[915] <= 0;
    valid_1[916]  <=   0;valid_2[916]  <=   0;dirty_bit_1[916] <= 0;dirty_bit_2[916] <= 0;lru_counter_1[916] <= 0;lru_counter_2[916] <= 0;tag_1[916] <= 0;tag_2[916] <= 0;cache_mem_1[916] <= 0;cache_mem_2[916] <= 0;
    valid_1[917]  <=   0;valid_2[917]  <=   0;dirty_bit_1[917] <= 0;dirty_bit_2[917] <= 0;lru_counter_1[917] <= 0;lru_counter_2[917] <= 0;tag_1[917] <= 0;tag_2[917] <= 0;cache_mem_1[917] <= 0;cache_mem_2[917] <= 0;
    valid_1[918]  <=   0;valid_2[918]  <=   0;dirty_bit_1[918] <= 0;dirty_bit_2[918] <= 0;lru_counter_1[918] <= 0;lru_counter_2[918] <= 0;tag_1[918] <= 0;tag_2[918] <= 0;cache_mem_1[918] <= 0;cache_mem_2[918] <= 0;
    valid_1[919]  <=   0;valid_2[919]  <=   0;dirty_bit_1[919] <= 0;dirty_bit_2[919] <= 0;lru_counter_1[919] <= 0;lru_counter_2[919] <= 0;tag_1[919] <= 0;tag_2[919] <= 0;cache_mem_1[919] <= 0;cache_mem_2[919] <= 0;
    valid_1[920]  <=   0;valid_2[920]  <=   0;dirty_bit_1[920] <= 0;dirty_bit_2[920] <= 0;lru_counter_1[920] <= 0;lru_counter_2[920] <= 0;tag_1[920] <= 0;tag_2[920] <= 0;cache_mem_1[920] <= 0;cache_mem_2[920] <= 0;
    valid_1[921]  <=   0;valid_2[921]  <=   0;dirty_bit_1[921] <= 0;dirty_bit_2[921] <= 0;lru_counter_1[921] <= 0;lru_counter_2[921] <= 0;tag_1[921] <= 0;tag_2[921] <= 0;cache_mem_1[921] <= 0;cache_mem_2[921] <= 0;
    valid_1[922]  <=   0;valid_2[922]  <=   0;dirty_bit_1[922] <= 0;dirty_bit_2[922] <= 0;lru_counter_1[922] <= 0;lru_counter_2[922] <= 0;tag_1[922] <= 0;tag_2[922] <= 0;cache_mem_1[922] <= 0;cache_mem_2[922] <= 0;
    valid_1[923]  <=   0;valid_2[923]  <=   0;dirty_bit_1[923] <= 0;dirty_bit_2[923] <= 0;lru_counter_1[923] <= 0;lru_counter_2[923] <= 0;tag_1[923] <= 0;tag_2[923] <= 0;cache_mem_1[923] <= 0;cache_mem_2[923] <= 0;
    valid_1[924]  <=   0;valid_2[924]  <=   0;dirty_bit_1[924] <= 0;dirty_bit_2[924] <= 0;lru_counter_1[924] <= 0;lru_counter_2[924] <= 0;tag_1[924] <= 0;tag_2[924] <= 0;cache_mem_1[924] <= 0;cache_mem_2[924] <= 0;
    valid_1[925]  <=   0;valid_2[925]  <=   0;dirty_bit_1[925] <= 0;dirty_bit_2[925] <= 0;lru_counter_1[925] <= 0;lru_counter_2[925] <= 0;tag_1[925] <= 0;tag_2[925] <= 0;cache_mem_1[925] <= 0;cache_mem_2[925] <= 0;
    valid_1[926]  <=   0;valid_2[926]  <=   0;dirty_bit_1[926] <= 0;dirty_bit_2[926] <= 0;lru_counter_1[926] <= 0;lru_counter_2[926] <= 0;tag_1[926] <= 0;tag_2[926] <= 0;cache_mem_1[926] <= 0;cache_mem_2[926] <= 0;
    valid_1[927]  <=   0;valid_2[927]  <=   0;dirty_bit_1[927] <= 0;dirty_bit_2[927] <= 0;lru_counter_1[927] <= 0;lru_counter_2[927] <= 0;tag_1[927] <= 0;tag_2[927] <= 0;cache_mem_1[927] <= 0;cache_mem_2[927] <= 0;
    valid_1[928]  <=   0;valid_2[928]  <=   0;dirty_bit_1[928] <= 0;dirty_bit_2[928] <= 0;lru_counter_1[928] <= 0;lru_counter_2[928] <= 0;tag_1[928] <= 0;tag_2[928] <= 0;cache_mem_1[928] <= 0;cache_mem_2[928] <= 0;
    valid_1[929]  <=   0;valid_2[929]  <=   0;dirty_bit_1[929] <= 0;dirty_bit_2[929] <= 0;lru_counter_1[929] <= 0;lru_counter_2[929] <= 0;tag_1[929] <= 0;tag_2[929] <= 0;cache_mem_1[929] <= 0;cache_mem_2[929] <= 0;
    valid_1[930]  <=   0;valid_2[930]  <=   0;dirty_bit_1[930] <= 0;dirty_bit_2[930] <= 0;lru_counter_1[930] <= 0;lru_counter_2[930] <= 0;tag_1[930] <= 0;tag_2[930] <= 0;cache_mem_1[930] <= 0;cache_mem_2[930] <= 0;
    valid_1[931]  <=   0;valid_2[931]  <=   0;dirty_bit_1[931] <= 0;dirty_bit_2[931] <= 0;lru_counter_1[931] <= 0;lru_counter_2[931] <= 0;tag_1[931] <= 0;tag_2[931] <= 0;cache_mem_1[931] <= 0;cache_mem_2[931] <= 0;
    valid_1[932]  <=   0;valid_2[932]  <=   0;dirty_bit_1[932] <= 0;dirty_bit_2[932] <= 0;lru_counter_1[932] <= 0;lru_counter_2[932] <= 0;tag_1[932] <= 0;tag_2[932] <= 0;cache_mem_1[932] <= 0;cache_mem_2[932] <= 0;
    valid_1[933]  <=   0;valid_2[933]  <=   0;dirty_bit_1[933] <= 0;dirty_bit_2[933] <= 0;lru_counter_1[933] <= 0;lru_counter_2[933] <= 0;tag_1[933] <= 0;tag_2[933] <= 0;cache_mem_1[933] <= 0;cache_mem_2[933] <= 0;
    valid_1[934]  <=   0;valid_2[934]  <=   0;dirty_bit_1[934] <= 0;dirty_bit_2[934] <= 0;lru_counter_1[934] <= 0;lru_counter_2[934] <= 0;tag_1[934] <= 0;tag_2[934] <= 0;cache_mem_1[934] <= 0;cache_mem_2[934] <= 0;
    valid_1[935]  <=   0;valid_2[935]  <=   0;dirty_bit_1[935] <= 0;dirty_bit_2[935] <= 0;lru_counter_1[935] <= 0;lru_counter_2[935] <= 0;tag_1[935] <= 0;tag_2[935] <= 0;cache_mem_1[935] <= 0;cache_mem_2[935] <= 0;
    valid_1[936]  <=   0;valid_2[936]  <=   0;dirty_bit_1[936] <= 0;dirty_bit_2[936] <= 0;lru_counter_1[936] <= 0;lru_counter_2[936] <= 0;tag_1[936] <= 0;tag_2[936] <= 0;cache_mem_1[936] <= 0;cache_mem_2[936] <= 0;
    valid_1[937]  <=   0;valid_2[937]  <=   0;dirty_bit_1[937] <= 0;dirty_bit_2[937] <= 0;lru_counter_1[937] <= 0;lru_counter_2[937] <= 0;tag_1[937] <= 0;tag_2[937] <= 0;cache_mem_1[937] <= 0;cache_mem_2[937] <= 0;
    valid_1[938]  <=   0;valid_2[938]  <=   0;dirty_bit_1[938] <= 0;dirty_bit_2[938] <= 0;lru_counter_1[938] <= 0;lru_counter_2[938] <= 0;tag_1[938] <= 0;tag_2[938] <= 0;cache_mem_1[938] <= 0;cache_mem_2[938] <= 0;
    valid_1[939]  <=   0;valid_2[939]  <=   0;dirty_bit_1[939] <= 0;dirty_bit_2[939] <= 0;lru_counter_1[939] <= 0;lru_counter_2[939] <= 0;tag_1[939] <= 0;tag_2[939] <= 0;cache_mem_1[939] <= 0;cache_mem_2[939] <= 0;
    valid_1[940]  <=   0;valid_2[940]  <=   0;dirty_bit_1[940] <= 0;dirty_bit_2[940] <= 0;lru_counter_1[940] <= 0;lru_counter_2[940] <= 0;tag_1[940] <= 0;tag_2[940] <= 0;cache_mem_1[940] <= 0;cache_mem_2[940] <= 0;
    valid_1[941]  <=   0;valid_2[941]  <=   0;dirty_bit_1[941] <= 0;dirty_bit_2[941] <= 0;lru_counter_1[941] <= 0;lru_counter_2[941] <= 0;tag_1[941] <= 0;tag_2[941] <= 0;cache_mem_1[941] <= 0;cache_mem_2[941] <= 0;
    valid_1[942]  <=   0;valid_2[942]  <=   0;dirty_bit_1[942] <= 0;dirty_bit_2[942] <= 0;lru_counter_1[942] <= 0;lru_counter_2[942] <= 0;tag_1[942] <= 0;tag_2[942] <= 0;cache_mem_1[942] <= 0;cache_mem_2[942] <= 0;
    valid_1[943]  <=   0;valid_2[943]  <=   0;dirty_bit_1[943] <= 0;dirty_bit_2[943] <= 0;lru_counter_1[943] <= 0;lru_counter_2[943] <= 0;tag_1[943] <= 0;tag_2[943] <= 0;cache_mem_1[943] <= 0;cache_mem_2[943] <= 0;
    valid_1[944]  <=   0;valid_2[944]  <=   0;dirty_bit_1[944] <= 0;dirty_bit_2[944] <= 0;lru_counter_1[944] <= 0;lru_counter_2[944] <= 0;tag_1[944] <= 0;tag_2[944] <= 0;cache_mem_1[944] <= 0;cache_mem_2[944] <= 0;
    valid_1[945]  <=   0;valid_2[945]  <=   0;dirty_bit_1[945] <= 0;dirty_bit_2[945] <= 0;lru_counter_1[945] <= 0;lru_counter_2[945] <= 0;tag_1[945] <= 0;tag_2[945] <= 0;cache_mem_1[945] <= 0;cache_mem_2[945] <= 0;
    valid_1[946]  <=   0;valid_2[946]  <=   0;dirty_bit_1[946] <= 0;dirty_bit_2[946] <= 0;lru_counter_1[946] <= 0;lru_counter_2[946] <= 0;tag_1[946] <= 0;tag_2[946] <= 0;cache_mem_1[946] <= 0;cache_mem_2[946] <= 0;
    valid_1[947]  <=   0;valid_2[947]  <=   0;dirty_bit_1[947] <= 0;dirty_bit_2[947] <= 0;lru_counter_1[947] <= 0;lru_counter_2[947] <= 0;tag_1[947] <= 0;tag_2[947] <= 0;cache_mem_1[947] <= 0;cache_mem_2[947] <= 0;
    valid_1[948]  <=   0;valid_2[948]  <=   0;dirty_bit_1[948] <= 0;dirty_bit_2[948] <= 0;lru_counter_1[948] <= 0;lru_counter_2[948] <= 0;tag_1[948] <= 0;tag_2[948] <= 0;cache_mem_1[948] <= 0;cache_mem_2[948] <= 0;
    valid_1[949]  <=   0;valid_2[949]  <=   0;dirty_bit_1[949] <= 0;dirty_bit_2[949] <= 0;lru_counter_1[949] <= 0;lru_counter_2[949] <= 0;tag_1[949] <= 0;tag_2[949] <= 0;cache_mem_1[949] <= 0;cache_mem_2[949] <= 0;
    valid_1[950]  <=   0;valid_2[950]  <=   0;dirty_bit_1[950] <= 0;dirty_bit_2[950] <= 0;lru_counter_1[950] <= 0;lru_counter_2[950] <= 0;tag_1[950] <= 0;tag_2[950] <= 0;cache_mem_1[950] <= 0;cache_mem_2[950] <= 0;
    valid_1[951]  <=   0;valid_2[951]  <=   0;dirty_bit_1[951] <= 0;dirty_bit_2[951] <= 0;lru_counter_1[951] <= 0;lru_counter_2[951] <= 0;tag_1[951] <= 0;tag_2[951] <= 0;cache_mem_1[951] <= 0;cache_mem_2[951] <= 0;
    valid_1[952]  <=   0;valid_2[952]  <=   0;dirty_bit_1[952] <= 0;dirty_bit_2[952] <= 0;lru_counter_1[952] <= 0;lru_counter_2[952] <= 0;tag_1[952] <= 0;tag_2[952] <= 0;cache_mem_1[952] <= 0;cache_mem_2[952] <= 0;
    valid_1[953]  <=   0;valid_2[953]  <=   0;dirty_bit_1[953] <= 0;dirty_bit_2[953] <= 0;lru_counter_1[953] <= 0;lru_counter_2[953] <= 0;tag_1[953] <= 0;tag_2[953] <= 0;cache_mem_1[953] <= 0;cache_mem_2[953] <= 0;
    valid_1[954]  <=   0;valid_2[954]  <=   0;dirty_bit_1[954] <= 0;dirty_bit_2[954] <= 0;lru_counter_1[954] <= 0;lru_counter_2[954] <= 0;tag_1[954] <= 0;tag_2[954] <= 0;cache_mem_1[954] <= 0;cache_mem_2[954] <= 0;
    valid_1[955]  <=   0;valid_2[955]  <=   0;dirty_bit_1[955] <= 0;dirty_bit_2[955] <= 0;lru_counter_1[955] <= 0;lru_counter_2[955] <= 0;tag_1[955] <= 0;tag_2[955] <= 0;cache_mem_1[955] <= 0;cache_mem_2[955] <= 0;
    valid_1[956]  <=   0;valid_2[956]  <=   0;dirty_bit_1[956] <= 0;dirty_bit_2[956] <= 0;lru_counter_1[956] <= 0;lru_counter_2[956] <= 0;tag_1[956] <= 0;tag_2[956] <= 0;cache_mem_1[956] <= 0;cache_mem_2[956] <= 0;
    valid_1[957]  <=   0;valid_2[957]  <=   0;dirty_bit_1[957] <= 0;dirty_bit_2[957] <= 0;lru_counter_1[957] <= 0;lru_counter_2[957] <= 0;tag_1[957] <= 0;tag_2[957] <= 0;cache_mem_1[957] <= 0;cache_mem_2[957] <= 0;
    valid_1[958]  <=   0;valid_2[958]  <=   0;dirty_bit_1[958] <= 0;dirty_bit_2[958] <= 0;lru_counter_1[958] <= 0;lru_counter_2[958] <= 0;tag_1[958] <= 0;tag_2[958] <= 0;cache_mem_1[958] <= 0;cache_mem_2[958] <= 0;
    valid_1[959]  <=   0;valid_2[959]  <=   0;dirty_bit_1[959] <= 0;dirty_bit_2[959] <= 0;lru_counter_1[959] <= 0;lru_counter_2[959] <= 0;tag_1[959] <= 0;tag_2[959] <= 0;cache_mem_1[959] <= 0;cache_mem_2[959] <= 0;
    valid_1[960]  <=   0;valid_2[960]  <=   0;dirty_bit_1[960] <= 0;dirty_bit_2[960] <= 0;lru_counter_1[960] <= 0;lru_counter_2[960] <= 0;tag_1[960] <= 0;tag_2[960] <= 0;cache_mem_1[960] <= 0;cache_mem_2[960] <= 0;
    valid_1[961]  <=   0;valid_2[961]  <=   0;dirty_bit_1[961] <= 0;dirty_bit_2[961] <= 0;lru_counter_1[961] <= 0;lru_counter_2[961] <= 0;tag_1[961] <= 0;tag_2[961] <= 0;cache_mem_1[961] <= 0;cache_mem_2[961] <= 0;
    valid_1[962]  <=   0;valid_2[962]  <=   0;dirty_bit_1[962] <= 0;dirty_bit_2[962] <= 0;lru_counter_1[962] <= 0;lru_counter_2[962] <= 0;tag_1[962] <= 0;tag_2[962] <= 0;cache_mem_1[962] <= 0;cache_mem_2[962] <= 0;
    valid_1[963]  <=   0;valid_2[963]  <=   0;dirty_bit_1[963] <= 0;dirty_bit_2[963] <= 0;lru_counter_1[963] <= 0;lru_counter_2[963] <= 0;tag_1[963] <= 0;tag_2[963] <= 0;cache_mem_1[963] <= 0;cache_mem_2[963] <= 0;
    valid_1[964]  <=   0;valid_2[964]  <=   0;dirty_bit_1[964] <= 0;dirty_bit_2[964] <= 0;lru_counter_1[964] <= 0;lru_counter_2[964] <= 0;tag_1[964] <= 0;tag_2[964] <= 0;cache_mem_1[964] <= 0;cache_mem_2[964] <= 0;
    valid_1[965]  <=   0;valid_2[965]  <=   0;dirty_bit_1[965] <= 0;dirty_bit_2[965] <= 0;lru_counter_1[965] <= 0;lru_counter_2[965] <= 0;tag_1[965] <= 0;tag_2[965] <= 0;cache_mem_1[965] <= 0;cache_mem_2[965] <= 0;
    valid_1[966]  <=   0;valid_2[966]  <=   0;dirty_bit_1[966] <= 0;dirty_bit_2[966] <= 0;lru_counter_1[966] <= 0;lru_counter_2[966] <= 0;tag_1[966] <= 0;tag_2[966] <= 0;cache_mem_1[966] <= 0;cache_mem_2[966] <= 0;
    valid_1[967]  <=   0;valid_2[967]  <=   0;dirty_bit_1[967] <= 0;dirty_bit_2[967] <= 0;lru_counter_1[967] <= 0;lru_counter_2[967] <= 0;tag_1[967] <= 0;tag_2[967] <= 0;cache_mem_1[967] <= 0;cache_mem_2[967] <= 0;
    valid_1[968]  <=   0;valid_2[968]  <=   0;dirty_bit_1[968] <= 0;dirty_bit_2[968] <= 0;lru_counter_1[968] <= 0;lru_counter_2[968] <= 0;tag_1[968] <= 0;tag_2[968] <= 0;cache_mem_1[968] <= 0;cache_mem_2[968] <= 0;
    valid_1[969]  <=   0;valid_2[969]  <=   0;dirty_bit_1[969] <= 0;dirty_bit_2[969] <= 0;lru_counter_1[969] <= 0;lru_counter_2[969] <= 0;tag_1[969] <= 0;tag_2[969] <= 0;cache_mem_1[969] <= 0;cache_mem_2[969] <= 0;
    valid_1[970]  <=   0;valid_2[970]  <=   0;dirty_bit_1[970] <= 0;dirty_bit_2[970] <= 0;lru_counter_1[970] <= 0;lru_counter_2[970] <= 0;tag_1[970] <= 0;tag_2[970] <= 0;cache_mem_1[970] <= 0;cache_mem_2[970] <= 0;
    valid_1[971]  <=   0;valid_2[971]  <=   0;dirty_bit_1[971] <= 0;dirty_bit_2[971] <= 0;lru_counter_1[971] <= 0;lru_counter_2[971] <= 0;tag_1[971] <= 0;tag_2[971] <= 0;cache_mem_1[971] <= 0;cache_mem_2[971] <= 0;
    valid_1[972]  <=   0;valid_2[972]  <=   0;dirty_bit_1[972] <= 0;dirty_bit_2[972] <= 0;lru_counter_1[972] <= 0;lru_counter_2[972] <= 0;tag_1[972] <= 0;tag_2[972] <= 0;cache_mem_1[972] <= 0;cache_mem_2[972] <= 0;
    valid_1[973]  <=   0;valid_2[973]  <=   0;dirty_bit_1[973] <= 0;dirty_bit_2[973] <= 0;lru_counter_1[973] <= 0;lru_counter_2[973] <= 0;tag_1[973] <= 0;tag_2[973] <= 0;cache_mem_1[973] <= 0;cache_mem_2[973] <= 0;
    valid_1[974]  <=   0;valid_2[974]  <=   0;dirty_bit_1[974] <= 0;dirty_bit_2[974] <= 0;lru_counter_1[974] <= 0;lru_counter_2[974] <= 0;tag_1[974] <= 0;tag_2[974] <= 0;cache_mem_1[974] <= 0;cache_mem_2[974] <= 0;
    valid_1[975]  <=   0;valid_2[975]  <=   0;dirty_bit_1[975] <= 0;dirty_bit_2[975] <= 0;lru_counter_1[975] <= 0;lru_counter_2[975] <= 0;tag_1[975] <= 0;tag_2[975] <= 0;cache_mem_1[975] <= 0;cache_mem_2[975] <= 0;
    valid_1[976]  <=   0;valid_2[976]  <=   0;dirty_bit_1[976] <= 0;dirty_bit_2[976] <= 0;lru_counter_1[976] <= 0;lru_counter_2[976] <= 0;tag_1[976] <= 0;tag_2[976] <= 0;cache_mem_1[976] <= 0;cache_mem_2[976] <= 0;
    valid_1[977]  <=   0;valid_2[977]  <=   0;dirty_bit_1[977] <= 0;dirty_bit_2[977] <= 0;lru_counter_1[977] <= 0;lru_counter_2[977] <= 0;tag_1[977] <= 0;tag_2[977] <= 0;cache_mem_1[977] <= 0;cache_mem_2[977] <= 0;
    valid_1[978]  <=   0;valid_2[978]  <=   0;dirty_bit_1[978] <= 0;dirty_bit_2[978] <= 0;lru_counter_1[978] <= 0;lru_counter_2[978] <= 0;tag_1[978] <= 0;tag_2[978] <= 0;cache_mem_1[978] <= 0;cache_mem_2[978] <= 0;
    valid_1[979]  <=   0;valid_2[979]  <=   0;dirty_bit_1[979] <= 0;dirty_bit_2[979] <= 0;lru_counter_1[979] <= 0;lru_counter_2[979] <= 0;tag_1[979] <= 0;tag_2[979] <= 0;cache_mem_1[979] <= 0;cache_mem_2[979] <= 0;
    valid_1[980]  <=   0;valid_2[980]  <=   0;dirty_bit_1[980] <= 0;dirty_bit_2[980] <= 0;lru_counter_1[980] <= 0;lru_counter_2[980] <= 0;tag_1[980] <= 0;tag_2[980] <= 0;cache_mem_1[980] <= 0;cache_mem_2[980] <= 0;
    valid_1[981]  <=   0;valid_2[981]  <=   0;dirty_bit_1[981] <= 0;dirty_bit_2[981] <= 0;lru_counter_1[981] <= 0;lru_counter_2[981] <= 0;tag_1[981] <= 0;tag_2[981] <= 0;cache_mem_1[981] <= 0;cache_mem_2[981] <= 0;
    valid_1[982]  <=   0;valid_2[982]  <=   0;dirty_bit_1[982] <= 0;dirty_bit_2[982] <= 0;lru_counter_1[982] <= 0;lru_counter_2[982] <= 0;tag_1[982] <= 0;tag_2[982] <= 0;cache_mem_1[982] <= 0;cache_mem_2[982] <= 0;
    valid_1[983]  <=   0;valid_2[983]  <=   0;dirty_bit_1[983] <= 0;dirty_bit_2[983] <= 0;lru_counter_1[983] <= 0;lru_counter_2[983] <= 0;tag_1[983] <= 0;tag_2[983] <= 0;cache_mem_1[983] <= 0;cache_mem_2[983] <= 0;
    valid_1[984]  <=   0;valid_2[984]  <=   0;dirty_bit_1[984] <= 0;dirty_bit_2[984] <= 0;lru_counter_1[984] <= 0;lru_counter_2[984] <= 0;tag_1[984] <= 0;tag_2[984] <= 0;cache_mem_1[984] <= 0;cache_mem_2[984] <= 0;
    valid_1[985]  <=   0;valid_2[985]  <=   0;dirty_bit_1[985] <= 0;dirty_bit_2[985] <= 0;lru_counter_1[985] <= 0;lru_counter_2[985] <= 0;tag_1[985] <= 0;tag_2[985] <= 0;cache_mem_1[985] <= 0;cache_mem_2[985] <= 0;
    valid_1[986]  <=   0;valid_2[986]  <=   0;dirty_bit_1[986] <= 0;dirty_bit_2[986] <= 0;lru_counter_1[986] <= 0;lru_counter_2[986] <= 0;tag_1[986] <= 0;tag_2[986] <= 0;cache_mem_1[986] <= 0;cache_mem_2[986] <= 0;
    valid_1[987]  <=   0;valid_2[987]  <=   0;dirty_bit_1[987] <= 0;dirty_bit_2[987] <= 0;lru_counter_1[987] <= 0;lru_counter_2[987] <= 0;tag_1[987] <= 0;tag_2[987] <= 0;cache_mem_1[987] <= 0;cache_mem_2[987] <= 0;
    valid_1[988]  <=   0;valid_2[988]  <=   0;dirty_bit_1[988] <= 0;dirty_bit_2[988] <= 0;lru_counter_1[988] <= 0;lru_counter_2[988] <= 0;tag_1[988] <= 0;tag_2[988] <= 0;cache_mem_1[988] <= 0;cache_mem_2[988] <= 0;
    valid_1[989]  <=   0;valid_2[989]  <=   0;dirty_bit_1[989] <= 0;dirty_bit_2[989] <= 0;lru_counter_1[989] <= 0;lru_counter_2[989] <= 0;tag_1[989] <= 0;tag_2[989] <= 0;cache_mem_1[989] <= 0;cache_mem_2[989] <= 0;
    valid_1[990]  <=   0;valid_2[990]  <=   0;dirty_bit_1[990] <= 0;dirty_bit_2[990] <= 0;lru_counter_1[990] <= 0;lru_counter_2[990] <= 0;tag_1[990] <= 0;tag_2[990] <= 0;cache_mem_1[990] <= 0;cache_mem_2[990] <= 0;
    valid_1[991]  <=   0;valid_2[991]  <=   0;dirty_bit_1[991] <= 0;dirty_bit_2[991] <= 0;lru_counter_1[991] <= 0;lru_counter_2[991] <= 0;tag_1[991] <= 0;tag_2[991] <= 0;cache_mem_1[991] <= 0;cache_mem_2[991] <= 0;
    valid_1[992]  <=   0;valid_2[992]  <=   0;dirty_bit_1[992] <= 0;dirty_bit_2[992] <= 0;lru_counter_1[992] <= 0;lru_counter_2[992] <= 0;tag_1[992] <= 0;tag_2[992] <= 0;cache_mem_1[992] <= 0;cache_mem_2[992] <= 0;
    valid_1[993]  <=   0;valid_2[993]  <=   0;dirty_bit_1[993] <= 0;dirty_bit_2[993] <= 0;lru_counter_1[993] <= 0;lru_counter_2[993] <= 0;tag_1[993] <= 0;tag_2[993] <= 0;cache_mem_1[993] <= 0;cache_mem_2[993] <= 0;
    valid_1[994]  <=   0;valid_2[994]  <=   0;dirty_bit_1[994] <= 0;dirty_bit_2[994] <= 0;lru_counter_1[994] <= 0;lru_counter_2[994] <= 0;tag_1[994] <= 0;tag_2[994] <= 0;cache_mem_1[994] <= 0;cache_mem_2[994] <= 0;
    valid_1[995]  <=   0;valid_2[995]  <=   0;dirty_bit_1[995] <= 0;dirty_bit_2[995] <= 0;lru_counter_1[995] <= 0;lru_counter_2[995] <= 0;tag_1[995] <= 0;tag_2[995] <= 0;cache_mem_1[995] <= 0;cache_mem_2[995] <= 0;
    valid_1[996]  <=   0;valid_2[996]  <=   0;dirty_bit_1[996] <= 0;dirty_bit_2[996] <= 0;lru_counter_1[996] <= 0;lru_counter_2[996] <= 0;tag_1[996] <= 0;tag_2[996] <= 0;cache_mem_1[996] <= 0;cache_mem_2[996] <= 0;
    valid_1[997]  <=   0;valid_2[997]  <=   0;dirty_bit_1[997] <= 0;dirty_bit_2[997] <= 0;lru_counter_1[997] <= 0;lru_counter_2[997] <= 0;tag_1[997] <= 0;tag_2[997] <= 0;cache_mem_1[997] <= 0;cache_mem_2[997] <= 0;
    valid_1[998]  <=   0;valid_2[998]  <=   0;dirty_bit_1[998] <= 0;dirty_bit_2[998] <= 0;lru_counter_1[998] <= 0;lru_counter_2[998] <= 0;tag_1[998] <= 0;tag_2[998] <= 0;cache_mem_1[998] <= 0;cache_mem_2[998] <= 0;
    valid_1[999]  <=   0;valid_2[999]  <=   0;dirty_bit_1[999] <= 0;dirty_bit_2[999] <= 0;lru_counter_1[999] <= 0;lru_counter_2[999] <= 0;tag_1[999] <= 0;tag_2[999] <= 0;cache_mem_1[999] <= 0;cache_mem_2[999] <= 0;
    valid_1[1000]  <=   0;valid_2[1000]  <=   0;dirty_bit_1[1000] <= 0;dirty_bit_2[1000] <= 0;lru_counter_1[1000] <= 0;lru_counter_2[1000] <= 0;tag_1[1000] <= 0;tag_2[1000] <= 0;cache_mem_1[1000] <= 0;cache_mem_2[1000] <= 0;
    valid_1[1001]  <=   0;valid_2[1001]  <=   0;dirty_bit_1[1001] <= 0;dirty_bit_2[1001] <= 0;lru_counter_1[1001] <= 0;lru_counter_2[1001] <= 0;tag_1[1001] <= 0;tag_2[1001] <= 0;cache_mem_1[1001] <= 0;cache_mem_2[1001] <= 0;
    valid_1[1002]  <=   0;valid_2[1002]  <=   0;dirty_bit_1[1002] <= 0;dirty_bit_2[1002] <= 0;lru_counter_1[1002] <= 0;lru_counter_2[1002] <= 0;tag_1[1002] <= 0;tag_2[1002] <= 0;cache_mem_1[1002] <= 0;cache_mem_2[1002] <= 0;
    valid_1[1003]  <=   0;valid_2[1003]  <=   0;dirty_bit_1[1003] <= 0;dirty_bit_2[1003] <= 0;lru_counter_1[1003] <= 0;lru_counter_2[1003] <= 0;tag_1[1003] <= 0;tag_2[1003] <= 0;cache_mem_1[1003] <= 0;cache_mem_2[1003] <= 0;
    valid_1[1004]  <=   0;valid_2[1004]  <=   0;dirty_bit_1[1004] <= 0;dirty_bit_2[1004] <= 0;lru_counter_1[1004] <= 0;lru_counter_2[1004] <= 0;tag_1[1004] <= 0;tag_2[1004] <= 0;cache_mem_1[1004] <= 0;cache_mem_2[1004] <= 0;
    valid_1[1005]  <=   0;valid_2[1005]  <=   0;dirty_bit_1[1005] <= 0;dirty_bit_2[1005] <= 0;lru_counter_1[1005] <= 0;lru_counter_2[1005] <= 0;tag_1[1005] <= 0;tag_2[1005] <= 0;cache_mem_1[1005] <= 0;cache_mem_2[1005] <= 0;
    valid_1[1006]  <=   0;valid_2[1006]  <=   0;dirty_bit_1[1006] <= 0;dirty_bit_2[1006] <= 0;lru_counter_1[1006] <= 0;lru_counter_2[1006] <= 0;tag_1[1006] <= 0;tag_2[1006] <= 0;cache_mem_1[1006] <= 0;cache_mem_2[1006] <= 0;
    valid_1[1007]  <=   0;valid_2[1007]  <=   0;dirty_bit_1[1007] <= 0;dirty_bit_2[1007] <= 0;lru_counter_1[1007] <= 0;lru_counter_2[1007] <= 0;tag_1[1007] <= 0;tag_2[1007] <= 0;cache_mem_1[1007] <= 0;cache_mem_2[1007] <= 0;
    valid_1[1008]  <=   0;valid_2[1008]  <=   0;dirty_bit_1[1008] <= 0;dirty_bit_2[1008] <= 0;lru_counter_1[1008] <= 0;lru_counter_2[1008] <= 0;tag_1[1008] <= 0;tag_2[1008] <= 0;cache_mem_1[1008] <= 0;cache_mem_2[1008] <= 0;
    valid_1[1009]  <=   0;valid_2[1009]  <=   0;dirty_bit_1[1009] <= 0;dirty_bit_2[1009] <= 0;lru_counter_1[1009] <= 0;lru_counter_2[1009] <= 0;tag_1[1009] <= 0;tag_2[1009] <= 0;cache_mem_1[1009] <= 0;cache_mem_2[1009] <= 0;
    valid_1[1010]  <=   0;valid_2[1010]  <=   0;dirty_bit_1[1010] <= 0;dirty_bit_2[1010] <= 0;lru_counter_1[1010] <= 0;lru_counter_2[1010] <= 0;tag_1[1010] <= 0;tag_2[1010] <= 0;cache_mem_1[1010] <= 0;cache_mem_2[1010] <= 0;
    valid_1[1011]  <=   0;valid_2[1011]  <=   0;dirty_bit_1[1011] <= 0;dirty_bit_2[1011] <= 0;lru_counter_1[1011] <= 0;lru_counter_2[1011] <= 0;tag_1[1011] <= 0;tag_2[1011] <= 0;cache_mem_1[1011] <= 0;cache_mem_2[1011] <= 0;
    valid_1[1012]  <=   0;valid_2[1012]  <=   0;dirty_bit_1[1012] <= 0;dirty_bit_2[1012] <= 0;lru_counter_1[1012] <= 0;lru_counter_2[1012] <= 0;tag_1[1012] <= 0;tag_2[1012] <= 0;cache_mem_1[1012] <= 0;cache_mem_2[1012] <= 0;
    valid_1[1013]  <=   0;valid_2[1013]  <=   0;dirty_bit_1[1013] <= 0;dirty_bit_2[1013] <= 0;lru_counter_1[1013] <= 0;lru_counter_2[1013] <= 0;tag_1[1013] <= 0;tag_2[1013] <= 0;cache_mem_1[1013] <= 0;cache_mem_2[1013] <= 0;
    valid_1[1014]  <=   0;valid_2[1014]  <=   0;dirty_bit_1[1014] <= 0;dirty_bit_2[1014] <= 0;lru_counter_1[1014] <= 0;lru_counter_2[1014] <= 0;tag_1[1014] <= 0;tag_2[1014] <= 0;cache_mem_1[1014] <= 0;cache_mem_2[1014] <= 0;
    valid_1[1015]  <=   0;valid_2[1015]  <=   0;dirty_bit_1[1015] <= 0;dirty_bit_2[1015] <= 0;lru_counter_1[1015] <= 0;lru_counter_2[1015] <= 0;tag_1[1015] <= 0;tag_2[1015] <= 0;cache_mem_1[1015] <= 0;cache_mem_2[1015] <= 0;
    valid_1[1016]  <=   0;valid_2[1016]  <=   0;dirty_bit_1[1016] <= 0;dirty_bit_2[1016] <= 0;lru_counter_1[1016] <= 0;lru_counter_2[1016] <= 0;tag_1[1016] <= 0;tag_2[1016] <= 0;cache_mem_1[1016] <= 0;cache_mem_2[1016] <= 0;
    valid_1[1017]  <=   0;valid_2[1017]  <=   0;dirty_bit_1[1017] <= 0;dirty_bit_2[1017] <= 0;lru_counter_1[1017] <= 0;lru_counter_2[1017] <= 0;tag_1[1017] <= 0;tag_2[1017] <= 0;cache_mem_1[1017] <= 0;cache_mem_2[1017] <= 0;
    valid_1[1018]  <=   0;valid_2[1018]  <=   0;dirty_bit_1[1018] <= 0;dirty_bit_2[1018] <= 0;lru_counter_1[1018] <= 0;lru_counter_2[1018] <= 0;tag_1[1018] <= 0;tag_2[1018] <= 0;cache_mem_1[1018] <= 0;cache_mem_2[1018] <= 0;
    valid_1[1019]  <=   0;valid_2[1019]  <=   0;dirty_bit_1[1019] <= 0;dirty_bit_2[1019] <= 0;lru_counter_1[1019] <= 0;lru_counter_2[1019] <= 0;tag_1[1019] <= 0;tag_2[1019] <= 0;cache_mem_1[1019] <= 0;cache_mem_2[1019] <= 0;
    valid_1[1020]  <=   0;valid_2[1020]  <=   0;dirty_bit_1[1020] <= 0;dirty_bit_2[1020] <= 0;lru_counter_1[1020] <= 0;lru_counter_2[1020] <= 0;tag_1[1020] <= 0;tag_2[1020] <= 0;cache_mem_1[1020] <= 0;cache_mem_2[1020] <= 0;
    valid_1[1021]  <=   0;valid_2[1021]  <=   0;dirty_bit_1[1021] <= 0;dirty_bit_2[1021] <= 0;lru_counter_1[1021] <= 0;lru_counter_2[1021] <= 0;tag_1[1021] <= 0;tag_2[1021] <= 0;cache_mem_1[1021] <= 0;cache_mem_2[1021] <= 0;
    valid_1[1022]  <=   0;valid_2[1022]  <=   0;dirty_bit_1[1022] <= 0;dirty_bit_2[1022] <= 0;lru_counter_1[1022] <= 0;lru_counter_2[1022] <= 0;tag_1[1022] <= 0;tag_2[1022] <= 0;cache_mem_1[1022] <= 0;cache_mem_2[1022] <= 0;
    valid_1[1023]  <=   0;valid_2[1023]  <=   0;dirty_bit_1[1023] <= 0;dirty_bit_2[1023] <= 0;lru_counter_1[1023] <= 0;lru_counter_2[1023] <= 0;tag_1[1023] <= 0;tag_2[1023] <= 0;cache_mem_1[1023] <= 0;cache_mem_2[1023] <= 0;
  end

end


endmodule



